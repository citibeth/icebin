netcdf _issm3 {
dimensions:
	grid.vertices.nrealized = 6708 ;
	grid.cells.nrealized = 12751 ;
	grid.cells.nrealized_plus1 = 12752 ;
	grid.cells.nvertex_refs = 38253 ;
	two = 2 ;
variables:
	int grid.info(two) ;
		grid.info:name = "ISSM_mesh" ;
		grid.info:version = 2 ;
		grid.info:type = "MESH" ;
		grid.info:coordinates = "XY" ;
		grid.info:parameterization = "L1" ;
		grid.info:projection = "+proj=stere +lon_0=-39 +lat_0=90 +lat_ts=71.0 +ellps=WGS84" ;
		grid.info:vertices.nfull = 6708 ;
		grid.info:cells.nfull = 12751 ;
	int grid.indexing(two) ;
		grid.indexing:base = 1 ;
		grid.indexing:extent = 6708 ;
		grid.indexing:indices = 0 ;
	int grid.vertices.index(grid.vertices.nrealized) ;
	double grid.vertices.xy(grid.vertices.nrealized, two) ;
	int grid.cells.index(grid.cells.nrealized) ;
	int grid.cells.vertex_refs(grid.cells.nvertex_refs) ;
	int grid.cells.vertex_refs_start(grid.cells.nrealized_plus1) ;
	double vertices.elevation(grid.vertices.nrealized) ;
data:

 grid.info = 
    1, 1 ;

 grid.indexing = 
    1, 1 ;

 grid.vertices.index = 
    1, 
    2, 
    3, 
    4, 
    5, 
    6, 
    7, 
    8, 
    9, 
    10, 
    11, 
    12, 
    13, 
    14, 
    15, 
    16, 
    17, 
    18, 
    19, 
    20, 
    21, 
    22, 
    23, 
    24, 
    25, 
    26, 
    27, 
    28, 
    29, 
    30, 
    31, 
    32, 
    33, 
    34, 
    35, 
    36, 
    37, 
    38, 
    39, 
    40, 
    41, 
    42, 
    43, 
    44, 
    45, 
    46, 
    47, 
    48, 
    49, 
    50, 
    51, 
    52, 
    53, 
    54, 
    55, 
    56, 
    57, 
    58, 
    59, 
    60, 
    61, 
    62, 
    63, 
    64, 
    65, 
    66, 
    67, 
    68, 
    69, 
    70, 
    71, 
    72, 
    73, 
    74, 
    75, 
    76, 
    77, 
    78, 
    79, 
    80, 
    81, 
    82, 
    83, 
    84, 
    85, 
    86, 
    87, 
    88, 
    89, 
    90, 
    91, 
    92, 
    93, 
    94, 
    95, 
    96, 
    97, 
    98, 
    99, 
    100, 
    101, 
    102, 
    103, 
    104, 
    105, 
    106, 
    107, 
    108, 
    109, 
    110, 
    111, 
    112, 
    113, 
    114, 
    115, 
    116, 
    117, 
    118, 
    119, 
    120, 
    121, 
    122, 
    123, 
    124, 
    125, 
    126, 
    127, 
    128, 
    129, 
    130, 
    131, 
    132, 
    133, 
    134, 
    135, 
    136, 
    137, 
    138, 
    139, 
    140, 
    141, 
    142, 
    143, 
    144, 
    145, 
    146, 
    147, 
    148, 
    149, 
    150, 
    151, 
    152, 
    153, 
    154, 
    155, 
    156, 
    157, 
    158, 
    159, 
    160, 
    161, 
    162, 
    163, 
    164, 
    165, 
    166, 
    167, 
    168, 
    169, 
    170, 
    171, 
    172, 
    173, 
    174, 
    175, 
    176, 
    177, 
    178, 
    179, 
    180, 
    181, 
    182, 
    183, 
    184, 
    185, 
    186, 
    187, 
    188, 
    189, 
    190, 
    191, 
    192, 
    193, 
    194, 
    195, 
    196, 
    197, 
    198, 
    199, 
    200, 
    201, 
    202, 
    203, 
    204, 
    205, 
    206, 
    207, 
    208, 
    209, 
    210, 
    211, 
    212, 
    213, 
    214, 
    215, 
    216, 
    217, 
    218, 
    219, 
    220, 
    221, 
    222, 
    223, 
    224, 
    225, 
    226, 
    227, 
    228, 
    229, 
    230, 
    231, 
    232, 
    233, 
    234, 
    235, 
    236, 
    237, 
    238, 
    239, 
    240, 
    241, 
    242, 
    243, 
    244, 
    245, 
    246, 
    247, 
    248, 
    249, 
    250, 
    251, 
    252, 
    253, 
    254, 
    255, 
    256, 
    257, 
    258, 
    259, 
    260, 
    261, 
    262, 
    263, 
    264, 
    265, 
    266, 
    267, 
    268, 
    269, 
    270, 
    271, 
    272, 
    273, 
    274, 
    275, 
    276, 
    277, 
    278, 
    279, 
    280, 
    281, 
    282, 
    283, 
    284, 
    285, 
    286, 
    287, 
    288, 
    289, 
    290, 
    291, 
    292, 
    293, 
    294, 
    295, 
    296, 
    297, 
    298, 
    299, 
    300, 
    301, 
    302, 
    303, 
    304, 
    305, 
    306, 
    307, 
    308, 
    309, 
    310, 
    311, 
    312, 
    313, 
    314, 
    315, 
    316, 
    317, 
    318, 
    319, 
    320, 
    321, 
    322, 
    323, 
    324, 
    325, 
    326, 
    327, 
    328, 
    329, 
    330, 
    331, 
    332, 
    333, 
    334, 
    335, 
    336, 
    337, 
    338, 
    339, 
    340, 
    341, 
    342, 
    343, 
    344, 
    345, 
    346, 
    347, 
    348, 
    349, 
    350, 
    351, 
    352, 
    353, 
    354, 
    355, 
    356, 
    357, 
    358, 
    359, 
    360, 
    361, 
    362, 
    363, 
    364, 
    365, 
    366, 
    367, 
    368, 
    369, 
    370, 
    371, 
    372, 
    373, 
    374, 
    375, 
    376, 
    377, 
    378, 
    379, 
    380, 
    381, 
    382, 
    383, 
    384, 
    385, 
    386, 
    387, 
    388, 
    389, 
    390, 
    391, 
    392, 
    393, 
    394, 
    395, 
    396, 
    397, 
    398, 
    399, 
    400, 
    401, 
    402, 
    403, 
    404, 
    405, 
    406, 
    407, 
    408, 
    409, 
    410, 
    411, 
    412, 
    413, 
    414, 
    415, 
    416, 
    417, 
    418, 
    419, 
    420, 
    421, 
    422, 
    423, 
    424, 
    425, 
    426, 
    427, 
    428, 
    429, 
    430, 
    431, 
    432, 
    433, 
    434, 
    435, 
    436, 
    437, 
    438, 
    439, 
    440, 
    441, 
    442, 
    443, 
    444, 
    445, 
    446, 
    447, 
    448, 
    449, 
    450, 
    451, 
    452, 
    453, 
    454, 
    455, 
    456, 
    457, 
    458, 
    459, 
    460, 
    461, 
    462, 
    463, 
    464, 
    465, 
    466, 
    467, 
    468, 
    469, 
    470, 
    471, 
    472, 
    473, 
    474, 
    475, 
    476, 
    477, 
    478, 
    479, 
    480, 
    481, 
    482, 
    483, 
    484, 
    485, 
    486, 
    487, 
    488, 
    489, 
    490, 
    491, 
    492, 
    493, 
    494, 
    495, 
    496, 
    497, 
    498, 
    499, 
    500, 
    501, 
    502, 
    503, 
    504, 
    505, 
    506, 
    507, 
    508, 
    509, 
    510, 
    511, 
    512, 
    513, 
    514, 
    515, 
    516, 
    517, 
    518, 
    519, 
    520, 
    521, 
    522, 
    523, 
    524, 
    525, 
    526, 
    527, 
    528, 
    529, 
    530, 
    531, 
    532, 
    533, 
    534, 
    535, 
    536, 
    537, 
    538, 
    539, 
    540, 
    541, 
    542, 
    543, 
    544, 
    545, 
    546, 
    547, 
    548, 
    549, 
    550, 
    551, 
    552, 
    553, 
    554, 
    555, 
    556, 
    557, 
    558, 
    559, 
    560, 
    561, 
    562, 
    563, 
    564, 
    565, 
    566, 
    567, 
    568, 
    569, 
    570, 
    571, 
    572, 
    573, 
    574, 
    575, 
    576, 
    577, 
    578, 
    579, 
    580, 
    581, 
    582, 
    583, 
    584, 
    585, 
    586, 
    587, 
    588, 
    589, 
    590, 
    591, 
    592, 
    593, 
    594, 
    595, 
    596, 
    597, 
    598, 
    599, 
    600, 
    601, 
    602, 
    603, 
    604, 
    605, 
    606, 
    607, 
    608, 
    609, 
    610, 
    611, 
    612, 
    613, 
    614, 
    615, 
    616, 
    617, 
    618, 
    619, 
    620, 
    621, 
    622, 
    623, 
    624, 
    625, 
    626, 
    627, 
    628, 
    629, 
    630, 
    631, 
    632, 
    633, 
    634, 
    635, 
    636, 
    637, 
    638, 
    639, 
    640, 
    641, 
    642, 
    643, 
    644, 
    645, 
    646, 
    647, 
    648, 
    649, 
    650, 
    651, 
    652, 
    653, 
    654, 
    655, 
    656, 
    657, 
    658, 
    659, 
    660, 
    661, 
    662, 
    663, 
    664, 
    665, 
    666, 
    667, 
    668, 
    669, 
    670, 
    671, 
    672, 
    673, 
    674, 
    675, 
    676, 
    677, 
    678, 
    679, 
    680, 
    681, 
    682, 
    683, 
    684, 
    685, 
    686, 
    687, 
    688, 
    689, 
    690, 
    691, 
    692, 
    693, 
    694, 
    695, 
    696, 
    697, 
    698, 
    699, 
    700, 
    701, 
    702, 
    703, 
    704, 
    705, 
    706, 
    707, 
    708, 
    709, 
    710, 
    711, 
    712, 
    713, 
    714, 
    715, 
    716, 
    717, 
    718, 
    719, 
    720, 
    721, 
    722, 
    723, 
    724, 
    725, 
    726, 
    727, 
    728, 
    729, 
    730, 
    731, 
    732, 
    733, 
    734, 
    735, 
    736, 
    737, 
    738, 
    739, 
    740, 
    741, 
    742, 
    743, 
    744, 
    745, 
    746, 
    747, 
    748, 
    749, 
    750, 
    751, 
    752, 
    753, 
    754, 
    755, 
    756, 
    757, 
    758, 
    759, 
    760, 
    761, 
    762, 
    763, 
    764, 
    765, 
    766, 
    767, 
    768, 
    769, 
    770, 
    771, 
    772, 
    773, 
    774, 
    775, 
    776, 
    777, 
    778, 
    779, 
    780, 
    781, 
    782, 
    783, 
    784, 
    785, 
    786, 
    787, 
    788, 
    789, 
    790, 
    791, 
    792, 
    793, 
    794, 
    795, 
    796, 
    797, 
    798, 
    799, 
    800, 
    801, 
    802, 
    803, 
    804, 
    805, 
    806, 
    807, 
    808, 
    809, 
    810, 
    811, 
    812, 
    813, 
    814, 
    815, 
    816, 
    817, 
    818, 
    819, 
    820, 
    821, 
    822, 
    823, 
    824, 
    825, 
    826, 
    827, 
    828, 
    829, 
    830, 
    831, 
    832, 
    833, 
    834, 
    835, 
    836, 
    837, 
    838, 
    839, 
    840, 
    841, 
    842, 
    843, 
    844, 
    845, 
    846, 
    847, 
    848, 
    849, 
    850, 
    851, 
    852, 
    853, 
    854, 
    855, 
    856, 
    857, 
    858, 
    859, 
    860, 
    861, 
    862, 
    863, 
    864, 
    865, 
    866, 
    867, 
    868, 
    869, 
    870, 
    871, 
    872, 
    873, 
    874, 
    875, 
    876, 
    877, 
    878, 
    879, 
    880, 
    881, 
    882, 
    883, 
    884, 
    885, 
    886, 
    887, 
    888, 
    889, 
    890, 
    891, 
    892, 
    893, 
    894, 
    895, 
    896, 
    897, 
    898, 
    899, 
    900, 
    901, 
    902, 
    903, 
    904, 
    905, 
    906, 
    907, 
    908, 
    909, 
    910, 
    911, 
    912, 
    913, 
    914, 
    915, 
    916, 
    917, 
    918, 
    919, 
    920, 
    921, 
    922, 
    923, 
    924, 
    925, 
    926, 
    927, 
    928, 
    929, 
    930, 
    931, 
    932, 
    933, 
    934, 
    935, 
    936, 
    937, 
    938, 
    939, 
    940, 
    941, 
    942, 
    943, 
    944, 
    945, 
    946, 
    947, 
    948, 
    949, 
    950, 
    951, 
    952, 
    953, 
    954, 
    955, 
    956, 
    957, 
    958, 
    959, 
    960, 
    961, 
    962, 
    963, 
    964, 
    965, 
    966, 
    967, 
    968, 
    969, 
    970, 
    971, 
    972, 
    973, 
    974, 
    975, 
    976, 
    977, 
    978, 
    979, 
    980, 
    981, 
    982, 
    983, 
    984, 
    985, 
    986, 
    987, 
    988, 
    989, 
    990, 
    991, 
    992, 
    993, 
    994, 
    995, 
    996, 
    997, 
    998, 
    999, 
    1000, 
    1001, 
    1002, 
    1003, 
    1004, 
    1005, 
    1006, 
    1007, 
    1008, 
    1009, 
    1010, 
    1011, 
    1012, 
    1013, 
    1014, 
    1015, 
    1016, 
    1017, 
    1018, 
    1019, 
    1020, 
    1021, 
    1022, 
    1023, 
    1024, 
    1025, 
    1026, 
    1027, 
    1028, 
    1029, 
    1030, 
    1031, 
    1032, 
    1033, 
    1034, 
    1035, 
    1036, 
    1037, 
    1038, 
    1039, 
    1040, 
    1041, 
    1042, 
    1043, 
    1044, 
    1045, 
    1046, 
    1047, 
    1048, 
    1049, 
    1050, 
    1051, 
    1052, 
    1053, 
    1054, 
    1055, 
    1056, 
    1057, 
    1058, 
    1059, 
    1060, 
    1061, 
    1062, 
    1063, 
    1064, 
    1065, 
    1066, 
    1067, 
    1068, 
    1069, 
    1070, 
    1071, 
    1072, 
    1073, 
    1074, 
    1075, 
    1076, 
    1077, 
    1078, 
    1079, 
    1080, 
    1081, 
    1082, 
    1083, 
    1084, 
    1085, 
    1086, 
    1087, 
    1088, 
    1089, 
    1090, 
    1091, 
    1092, 
    1093, 
    1094, 
    1095, 
    1096, 
    1097, 
    1098, 
    1099, 
    1100, 
    1101, 
    1102, 
    1103, 
    1104, 
    1105, 
    1106, 
    1107, 
    1108, 
    1109, 
    1110, 
    1111, 
    1112, 
    1113, 
    1114, 
    1115, 
    1116, 
    1117, 
    1118, 
    1119, 
    1120, 
    1121, 
    1122, 
    1123, 
    1124, 
    1125, 
    1126, 
    1127, 
    1128, 
    1129, 
    1130, 
    1131, 
    1132, 
    1133, 
    1134, 
    1135, 
    1136, 
    1137, 
    1138, 
    1139, 
    1140, 
    1141, 
    1142, 
    1143, 
    1144, 
    1145, 
    1146, 
    1147, 
    1148, 
    1149, 
    1150, 
    1151, 
    1152, 
    1153, 
    1154, 
    1155, 
    1156, 
    1157, 
    1158, 
    1159, 
    1160, 
    1161, 
    1162, 
    1163, 
    1164, 
    1165, 
    1166, 
    1167, 
    1168, 
    1169, 
    1170, 
    1171, 
    1172, 
    1173, 
    1174, 
    1175, 
    1176, 
    1177, 
    1178, 
    1179, 
    1180, 
    1181, 
    1182, 
    1183, 
    1184, 
    1185, 
    1186, 
    1187, 
    1188, 
    1189, 
    1190, 
    1191, 
    1192, 
    1193, 
    1194, 
    1195, 
    1196, 
    1197, 
    1198, 
    1199, 
    1200, 
    1201, 
    1202, 
    1203, 
    1204, 
    1205, 
    1206, 
    1207, 
    1208, 
    1209, 
    1210, 
    1211, 
    1212, 
    1213, 
    1214, 
    1215, 
    1216, 
    1217, 
    1218, 
    1219, 
    1220, 
    1221, 
    1222, 
    1223, 
    1224, 
    1225, 
    1226, 
    1227, 
    1228, 
    1229, 
    1230, 
    1231, 
    1232, 
    1233, 
    1234, 
    1235, 
    1236, 
    1237, 
    1238, 
    1239, 
    1240, 
    1241, 
    1242, 
    1243, 
    1244, 
    1245, 
    1246, 
    1247, 
    1248, 
    1249, 
    1250, 
    1251, 
    1252, 
    1253, 
    1254, 
    1255, 
    1256, 
    1257, 
    1258, 
    1259, 
    1260, 
    1261, 
    1262, 
    1263, 
    1264, 
    1265, 
    1266, 
    1267, 
    1268, 
    1269, 
    1270, 
    1271, 
    1272, 
    1273, 
    1274, 
    1275, 
    1276, 
    1277, 
    1278, 
    1279, 
    1280, 
    1281, 
    1282, 
    1283, 
    1284, 
    1285, 
    1286, 
    1287, 
    1288, 
    1289, 
    1290, 
    1291, 
    1292, 
    1293, 
    1294, 
    1295, 
    1296, 
    1297, 
    1298, 
    1299, 
    1300, 
    1301, 
    1302, 
    1303, 
    1304, 
    1305, 
    1306, 
    1307, 
    1308, 
    1309, 
    1310, 
    1311, 
    1312, 
    1313, 
    1314, 
    1315, 
    1316, 
    1317, 
    1318, 
    1319, 
    1320, 
    1321, 
    1322, 
    1323, 
    1324, 
    1325, 
    1326, 
    1327, 
    1328, 
    1329, 
    1330, 
    1331, 
    1332, 
    1333, 
    1334, 
    1335, 
    1336, 
    1337, 
    1338, 
    1339, 
    1340, 
    1341, 
    1342, 
    1343, 
    1344, 
    1345, 
    1346, 
    1347, 
    1348, 
    1349, 
    1350, 
    1351, 
    1352, 
    1353, 
    1354, 
    1355, 
    1356, 
    1357, 
    1358, 
    1359, 
    1360, 
    1361, 
    1362, 
    1363, 
    1364, 
    1365, 
    1366, 
    1367, 
    1368, 
    1369, 
    1370, 
    1371, 
    1372, 
    1373, 
    1374, 
    1375, 
    1376, 
    1377, 
    1378, 
    1379, 
    1380, 
    1381, 
    1382, 
    1383, 
    1384, 
    1385, 
    1386, 
    1387, 
    1388, 
    1389, 
    1390, 
    1391, 
    1392, 
    1393, 
    1394, 
    1395, 
    1396, 
    1397, 
    1398, 
    1399, 
    1400, 
    1401, 
    1402, 
    1403, 
    1404, 
    1405, 
    1406, 
    1407, 
    1408, 
    1409, 
    1410, 
    1411, 
    1412, 
    1413, 
    1414, 
    1415, 
    1416, 
    1417, 
    1418, 
    1419, 
    1420, 
    1421, 
    1422, 
    1423, 
    1424, 
    1425, 
    1426, 
    1427, 
    1428, 
    1429, 
    1430, 
    1431, 
    1432, 
    1433, 
    1434, 
    1435, 
    1436, 
    1437, 
    1438, 
    1439, 
    1440, 
    1441, 
    1442, 
    1443, 
    1444, 
    1445, 
    1446, 
    1447, 
    1448, 
    1449, 
    1450, 
    1451, 
    1452, 
    1453, 
    1454, 
    1455, 
    1456, 
    1457, 
    1458, 
    1459, 
    1460, 
    1461, 
    1462, 
    1463, 
    1464, 
    1465, 
    1466, 
    1467, 
    1468, 
    1469, 
    1470, 
    1471, 
    1472, 
    1473, 
    1474, 
    1475, 
    1476, 
    1477, 
    1478, 
    1479, 
    1480, 
    1481, 
    1482, 
    1483, 
    1484, 
    1485, 
    1486, 
    1487, 
    1488, 
    1489, 
    1490, 
    1491, 
    1492, 
    1493, 
    1494, 
    1495, 
    1496, 
    1497, 
    1498, 
    1499, 
    1500, 
    1501, 
    1502, 
    1503, 
    1504, 
    1505, 
    1506, 
    1507, 
    1508, 
    1509, 
    1510, 
    1511, 
    1512, 
    1513, 
    1514, 
    1515, 
    1516, 
    1517, 
    1518, 
    1519, 
    1520, 
    1521, 
    1522, 
    1523, 
    1524, 
    1525, 
    1526, 
    1527, 
    1528, 
    1529, 
    1530, 
    1531, 
    1532, 
    1533, 
    1534, 
    1535, 
    1536, 
    1537, 
    1538, 
    1539, 
    1540, 
    1541, 
    1542, 
    1543, 
    1544, 
    1545, 
    1546, 
    1547, 
    1548, 
    1549, 
    1550, 
    1551, 
    1552, 
    1553, 
    1554, 
    1555, 
    1556, 
    1557, 
    1558, 
    1559, 
    1560, 
    1561, 
    1562, 
    1563, 
    1564, 
    1565, 
    1566, 
    1567, 
    1568, 
    1569, 
    1570, 
    1571, 
    1572, 
    1573, 
    1574, 
    1575, 
    1576, 
    1577, 
    1578, 
    1579, 
    1580, 
    1581, 
    1582, 
    1583, 
    1584, 
    1585, 
    1586, 
    1587, 
    1588, 
    1589, 
    1590, 
    1591, 
    1592, 
    1593, 
    1594, 
    1595, 
    1596, 
    1597, 
    1598, 
    1599, 
    1600, 
    1601, 
    1602, 
    1603, 
    1604, 
    1605, 
    1606, 
    1607, 
    1608, 
    1609, 
    1610, 
    1611, 
    1612, 
    1613, 
    1614, 
    1615, 
    1616, 
    1617, 
    1618, 
    1619, 
    1620, 
    1621, 
    1622, 
    1623, 
    1624, 
    1625, 
    1626, 
    1627, 
    1628, 
    1629, 
    1630, 
    1631, 
    1632, 
    1633, 
    1634, 
    1635, 
    1636, 
    1637, 
    1638, 
    1639, 
    1640, 
    1641, 
    1642, 
    1643, 
    1644, 
    1645, 
    1646, 
    1647, 
    1648, 
    1649, 
    1650, 
    1651, 
    1652, 
    1653, 
    1654, 
    1655, 
    1656, 
    1657, 
    1658, 
    1659, 
    1660, 
    1661, 
    1662, 
    1663, 
    1664, 
    1665, 
    1666, 
    1667, 
    1668, 
    1669, 
    1670, 
    1671, 
    1672, 
    1673, 
    1674, 
    1675, 
    1676, 
    1677, 
    1678, 
    1679, 
    1680, 
    1681, 
    1682, 
    1683, 
    1684, 
    1685, 
    1686, 
    1687, 
    1688, 
    1689, 
    1690, 
    1691, 
    1692, 
    1693, 
    1694, 
    1695, 
    1696, 
    1697, 
    1698, 
    1699, 
    1700, 
    1701, 
    1702, 
    1703, 
    1704, 
    1705, 
    1706, 
    1707, 
    1708, 
    1709, 
    1710, 
    1711, 
    1712, 
    1713, 
    1714, 
    1715, 
    1716, 
    1717, 
    1718, 
    1719, 
    1720, 
    1721, 
    1722, 
    1723, 
    1724, 
    1725, 
    1726, 
    1727, 
    1728, 
    1729, 
    1730, 
    1731, 
    1732, 
    1733, 
    1734, 
    1735, 
    1736, 
    1737, 
    1738, 
    1739, 
    1740, 
    1741, 
    1742, 
    1743, 
    1744, 
    1745, 
    1746, 
    1747, 
    1748, 
    1749, 
    1750, 
    1751, 
    1752, 
    1753, 
    1754, 
    1755, 
    1756, 
    1757, 
    1758, 
    1759, 
    1760, 
    1761, 
    1762, 
    1763, 
    1764, 
    1765, 
    1766, 
    1767, 
    1768, 
    1769, 
    1770, 
    1771, 
    1772, 
    1773, 
    1774, 
    1775, 
    1776, 
    1777, 
    1778, 
    1779, 
    1780, 
    1781, 
    1782, 
    1783, 
    1784, 
    1785, 
    1786, 
    1787, 
    1788, 
    1789, 
    1790, 
    1791, 
    1792, 
    1793, 
    1794, 
    1795, 
    1796, 
    1797, 
    1798, 
    1799, 
    1800, 
    1801, 
    1802, 
    1803, 
    1804, 
    1805, 
    1806, 
    1807, 
    1808, 
    1809, 
    1810, 
    1811, 
    1812, 
    1813, 
    1814, 
    1815, 
    1816, 
    1817, 
    1818, 
    1819, 
    1820, 
    1821, 
    1822, 
    1823, 
    1824, 
    1825, 
    1826, 
    1827, 
    1828, 
    1829, 
    1830, 
    1831, 
    1832, 
    1833, 
    1834, 
    1835, 
    1836, 
    1837, 
    1838, 
    1839, 
    1840, 
    1841, 
    1842, 
    1843, 
    1844, 
    1845, 
    1846, 
    1847, 
    1848, 
    1849, 
    1850, 
    1851, 
    1852, 
    1853, 
    1854, 
    1855, 
    1856, 
    1857, 
    1858, 
    1859, 
    1860, 
    1861, 
    1862, 
    1863, 
    1864, 
    1865, 
    1866, 
    1867, 
    1868, 
    1869, 
    1870, 
    1871, 
    1872, 
    1873, 
    1874, 
    1875, 
    1876, 
    1877, 
    1878, 
    1879, 
    1880, 
    1881, 
    1882, 
    1883, 
    1884, 
    1885, 
    1886, 
    1887, 
    1888, 
    1889, 
    1890, 
    1891, 
    1892, 
    1893, 
    1894, 
    1895, 
    1896, 
    1897, 
    1898, 
    1899, 
    1900, 
    1901, 
    1902, 
    1903, 
    1904, 
    1905, 
    1906, 
    1907, 
    1908, 
    1909, 
    1910, 
    1911, 
    1912, 
    1913, 
    1914, 
    1915, 
    1916, 
    1917, 
    1918, 
    1919, 
    1920, 
    1921, 
    1922, 
    1923, 
    1924, 
    1925, 
    1926, 
    1927, 
    1928, 
    1929, 
    1930, 
    1931, 
    1932, 
    1933, 
    1934, 
    1935, 
    1936, 
    1937, 
    1938, 
    1939, 
    1940, 
    1941, 
    1942, 
    1943, 
    1944, 
    1945, 
    1946, 
    1947, 
    1948, 
    1949, 
    1950, 
    1951, 
    1952, 
    1953, 
    1954, 
    1955, 
    1956, 
    1957, 
    1958, 
    1959, 
    1960, 
    1961, 
    1962, 
    1963, 
    1964, 
    1965, 
    1966, 
    1967, 
    1968, 
    1969, 
    1970, 
    1971, 
    1972, 
    1973, 
    1974, 
    1975, 
    1976, 
    1977, 
    1978, 
    1979, 
    1980, 
    1981, 
    1982, 
    1983, 
    1984, 
    1985, 
    1986, 
    1987, 
    1988, 
    1989, 
    1990, 
    1991, 
    1992, 
    1993, 
    1994, 
    1995, 
    1996, 
    1997, 
    1998, 
    1999, 
    2000, 
    2001, 
    2002, 
    2003, 
    2004, 
    2005, 
    2006, 
    2007, 
    2008, 
    2009, 
    2010, 
    2011, 
    2012, 
    2013, 
    2014, 
    2015, 
    2016, 
    2017, 
    2018, 
    2019, 
    2020, 
    2021, 
    2022, 
    2023, 
    2024, 
    2025, 
    2026, 
    2027, 
    2028, 
    2029, 
    2030, 
    2031, 
    2032, 
    2033, 
    2034, 
    2035, 
    2036, 
    2037, 
    2038, 
    2039, 
    2040, 
    2041, 
    2042, 
    2043, 
    2044, 
    2045, 
    2046, 
    2047, 
    2048, 
    2049, 
    2050, 
    2051, 
    2052, 
    2053, 
    2054, 
    2055, 
    2056, 
    2057, 
    2058, 
    2059, 
    2060, 
    2061, 
    2062, 
    2063, 
    2064, 
    2065, 
    2066, 
    2067, 
    2068, 
    2069, 
    2070, 
    2071, 
    2072, 
    2073, 
    2074, 
    2075, 
    2076, 
    2077, 
    2078, 
    2079, 
    2080, 
    2081, 
    2082, 
    2083, 
    2084, 
    2085, 
    2086, 
    2087, 
    2088, 
    2089, 
    2090, 
    2091, 
    2092, 
    2093, 
    2094, 
    2095, 
    2096, 
    2097, 
    2098, 
    2099, 
    2100, 
    2101, 
    2102, 
    2103, 
    2104, 
    2105, 
    2106, 
    2107, 
    2108, 
    2109, 
    2110, 
    2111, 
    2112, 
    2113, 
    2114, 
    2115, 
    2116, 
    2117, 
    2118, 
    2119, 
    2120, 
    2121, 
    2122, 
    2123, 
    2124, 
    2125, 
    2126, 
    2127, 
    2128, 
    2129, 
    2130, 
    2131, 
    2132, 
    2133, 
    2134, 
    2135, 
    2136, 
    2137, 
    2138, 
    2139, 
    2140, 
    2141, 
    2142, 
    2143, 
    2144, 
    2145, 
    2146, 
    2147, 
    2148, 
    2149, 
    2150, 
    2151, 
    2152, 
    2153, 
    2154, 
    2155, 
    2156, 
    2157, 
    2158, 
    2159, 
    2160, 
    2161, 
    2162, 
    2163, 
    2164, 
    2165, 
    2166, 
    2167, 
    2168, 
    2169, 
    2170, 
    2171, 
    2172, 
    2173, 
    2174, 
    2175, 
    2176, 
    2177, 
    2178, 
    2179, 
    2180, 
    2181, 
    2182, 
    2183, 
    2184, 
    2185, 
    2186, 
    2187, 
    2188, 
    2189, 
    2190, 
    2191, 
    2192, 
    2193, 
    2194, 
    2195, 
    2196, 
    2197, 
    2198, 
    2199, 
    2200, 
    2201, 
    2202, 
    2203, 
    2204, 
    2205, 
    2206, 
    2207, 
    2208, 
    2209, 
    2210, 
    2211, 
    2212, 
    2213, 
    2214, 
    2215, 
    2216, 
    2217, 
    2218, 
    2219, 
    2220, 
    2221, 
    2222, 
    2223, 
    2224, 
    2225, 
    2226, 
    2227, 
    2228, 
    2229, 
    2230, 
    2231, 
    2232, 
    2233, 
    2234, 
    2235, 
    2236, 
    2237, 
    2238, 
    2239, 
    2240, 
    2241, 
    2242, 
    2243, 
    2244, 
    2245, 
    2246, 
    2247, 
    2248, 
    2249, 
    2250, 
    2251, 
    2252, 
    2253, 
    2254, 
    2255, 
    2256, 
    2257, 
    2258, 
    2259, 
    2260, 
    2261, 
    2262, 
    2263, 
    2264, 
    2265, 
    2266, 
    2267, 
    2268, 
    2269, 
    2270, 
    2271, 
    2272, 
    2273, 
    2274, 
    2275, 
    2276, 
    2277, 
    2278, 
    2279, 
    2280, 
    2281, 
    2282, 
    2283, 
    2284, 
    2285, 
    2286, 
    2287, 
    2288, 
    2289, 
    2290, 
    2291, 
    2292, 
    2293, 
    2294, 
    2295, 
    2296, 
    2297, 
    2298, 
    2299, 
    2300, 
    2301, 
    2302, 
    2303, 
    2304, 
    2305, 
    2306, 
    2307, 
    2308, 
    2309, 
    2310, 
    2311, 
    2312, 
    2313, 
    2314, 
    2315, 
    2316, 
    2317, 
    2318, 
    2319, 
    2320, 
    2321, 
    2322, 
    2323, 
    2324, 
    2325, 
    2326, 
    2327, 
    2328, 
    2329, 
    2330, 
    2331, 
    2332, 
    2333, 
    2334, 
    2335, 
    2336, 
    2337, 
    2338, 
    2339, 
    2340, 
    2341, 
    2342, 
    2343, 
    2344, 
    2345, 
    2346, 
    2347, 
    2348, 
    2349, 
    2350, 
    2351, 
    2352, 
    2353, 
    2354, 
    2355, 
    2356, 
    2357, 
    2358, 
    2359, 
    2360, 
    2361, 
    2362, 
    2363, 
    2364, 
    2365, 
    2366, 
    2367, 
    2368, 
    2369, 
    2370, 
    2371, 
    2372, 
    2373, 
    2374, 
    2375, 
    2376, 
    2377, 
    2378, 
    2379, 
    2380, 
    2381, 
    2382, 
    2383, 
    2384, 
    2385, 
    2386, 
    2387, 
    2388, 
    2389, 
    2390, 
    2391, 
    2392, 
    2393, 
    2394, 
    2395, 
    2396, 
    2397, 
    2398, 
    2399, 
    2400, 
    2401, 
    2402, 
    2403, 
    2404, 
    2405, 
    2406, 
    2407, 
    2408, 
    2409, 
    2410, 
    2411, 
    2412, 
    2413, 
    2414, 
    2415, 
    2416, 
    2417, 
    2418, 
    2419, 
    2420, 
    2421, 
    2422, 
    2423, 
    2424, 
    2425, 
    2426, 
    2427, 
    2428, 
    2429, 
    2430, 
    2431, 
    2432, 
    2433, 
    2434, 
    2435, 
    2436, 
    2437, 
    2438, 
    2439, 
    2440, 
    2441, 
    2442, 
    2443, 
    2444, 
    2445, 
    2446, 
    2447, 
    2448, 
    2449, 
    2450, 
    2451, 
    2452, 
    2453, 
    2454, 
    2455, 
    2456, 
    2457, 
    2458, 
    2459, 
    2460, 
    2461, 
    2462, 
    2463, 
    2464, 
    2465, 
    2466, 
    2467, 
    2468, 
    2469, 
    2470, 
    2471, 
    2472, 
    2473, 
    2474, 
    2475, 
    2476, 
    2477, 
    2478, 
    2479, 
    2480, 
    2481, 
    2482, 
    2483, 
    2484, 
    2485, 
    2486, 
    2487, 
    2488, 
    2489, 
    2490, 
    2491, 
    2492, 
    2493, 
    2494, 
    2495, 
    2496, 
    2497, 
    2498, 
    2499, 
    2500, 
    2501, 
    2502, 
    2503, 
    2504, 
    2505, 
    2506, 
    2507, 
    2508, 
    2509, 
    2510, 
    2511, 
    2512, 
    2513, 
    2514, 
    2515, 
    2516, 
    2517, 
    2518, 
    2519, 
    2520, 
    2521, 
    2522, 
    2523, 
    2524, 
    2525, 
    2526, 
    2527, 
    2528, 
    2529, 
    2530, 
    2531, 
    2532, 
    2533, 
    2534, 
    2535, 
    2536, 
    2537, 
    2538, 
    2539, 
    2540, 
    2541, 
    2542, 
    2543, 
    2544, 
    2545, 
    2546, 
    2547, 
    2548, 
    2549, 
    2550, 
    2551, 
    2552, 
    2553, 
    2554, 
    2555, 
    2556, 
    2557, 
    2558, 
    2559, 
    2560, 
    2561, 
    2562, 
    2563, 
    2564, 
    2565, 
    2566, 
    2567, 
    2568, 
    2569, 
    2570, 
    2571, 
    2572, 
    2573, 
    2574, 
    2575, 
    2576, 
    2577, 
    2578, 
    2579, 
    2580, 
    2581, 
    2582, 
    2583, 
    2584, 
    2585, 
    2586, 
    2587, 
    2588, 
    2589, 
    2590, 
    2591, 
    2592, 
    2593, 
    2594, 
    2595, 
    2596, 
    2597, 
    2598, 
    2599, 
    2600, 
    2601, 
    2602, 
    2603, 
    2604, 
    2605, 
    2606, 
    2607, 
    2608, 
    2609, 
    2610, 
    2611, 
    2612, 
    2613, 
    2614, 
    2615, 
    2616, 
    2617, 
    2618, 
    2619, 
    2620, 
    2621, 
    2622, 
    2623, 
    2624, 
    2625, 
    2626, 
    2627, 
    2628, 
    2629, 
    2630, 
    2631, 
    2632, 
    2633, 
    2634, 
    2635, 
    2636, 
    2637, 
    2638, 
    2639, 
    2640, 
    2641, 
    2642, 
    2643, 
    2644, 
    2645, 
    2646, 
    2647, 
    2648, 
    2649, 
    2650, 
    2651, 
    2652, 
    2653, 
    2654, 
    2655, 
    2656, 
    2657, 
    2658, 
    2659, 
    2660, 
    2661, 
    2662, 
    2663, 
    2664, 
    2665, 
    2666, 
    2667, 
    2668, 
    2669, 
    2670, 
    2671, 
    2672, 
    2673, 
    2674, 
    2675, 
    2676, 
    2677, 
    2678, 
    2679, 
    2680, 
    2681, 
    2682, 
    2683, 
    2684, 
    2685, 
    2686, 
    2687, 
    2688, 
    2689, 
    2690, 
    2691, 
    2692, 
    2693, 
    2694, 
    2695, 
    2696, 
    2697, 
    2698, 
    2699, 
    2700, 
    2701, 
    2702, 
    2703, 
    2704, 
    2705, 
    2706, 
    2707, 
    2708, 
    2709, 
    2710, 
    2711, 
    2712, 
    2713, 
    2714, 
    2715, 
    2716, 
    2717, 
    2718, 
    2719, 
    2720, 
    2721, 
    2722, 
    2723, 
    2724, 
    2725, 
    2726, 
    2727, 
    2728, 
    2729, 
    2730, 
    2731, 
    2732, 
    2733, 
    2734, 
    2735, 
    2736, 
    2737, 
    2738, 
    2739, 
    2740, 
    2741, 
    2742, 
    2743, 
    2744, 
    2745, 
    2746, 
    2747, 
    2748, 
    2749, 
    2750, 
    2751, 
    2752, 
    2753, 
    2754, 
    2755, 
    2756, 
    2757, 
    2758, 
    2759, 
    2760, 
    2761, 
    2762, 
    2763, 
    2764, 
    2765, 
    2766, 
    2767, 
    2768, 
    2769, 
    2770, 
    2771, 
    2772, 
    2773, 
    2774, 
    2775, 
    2776, 
    2777, 
    2778, 
    2779, 
    2780, 
    2781, 
    2782, 
    2783, 
    2784, 
    2785, 
    2786, 
    2787, 
    2788, 
    2789, 
    2790, 
    2791, 
    2792, 
    2793, 
    2794, 
    2795, 
    2796, 
    2797, 
    2798, 
    2799, 
    2800, 
    2801, 
    2802, 
    2803, 
    2804, 
    2805, 
    2806, 
    2807, 
    2808, 
    2809, 
    2810, 
    2811, 
    2812, 
    2813, 
    2814, 
    2815, 
    2816, 
    2817, 
    2818, 
    2819, 
    2820, 
    2821, 
    2822, 
    2823, 
    2824, 
    2825, 
    2826, 
    2827, 
    2828, 
    2829, 
    2830, 
    2831, 
    2832, 
    2833, 
    2834, 
    2835, 
    2836, 
    2837, 
    2838, 
    2839, 
    2840, 
    2841, 
    2842, 
    2843, 
    2844, 
    2845, 
    2846, 
    2847, 
    2848, 
    2849, 
    2850, 
    2851, 
    2852, 
    2853, 
    2854, 
    2855, 
    2856, 
    2857, 
    2858, 
    2859, 
    2860, 
    2861, 
    2862, 
    2863, 
    2864, 
    2865, 
    2866, 
    2867, 
    2868, 
    2869, 
    2870, 
    2871, 
    2872, 
    2873, 
    2874, 
    2875, 
    2876, 
    2877, 
    2878, 
    2879, 
    2880, 
    2881, 
    2882, 
    2883, 
    2884, 
    2885, 
    2886, 
    2887, 
    2888, 
    2889, 
    2890, 
    2891, 
    2892, 
    2893, 
    2894, 
    2895, 
    2896, 
    2897, 
    2898, 
    2899, 
    2900, 
    2901, 
    2902, 
    2903, 
    2904, 
    2905, 
    2906, 
    2907, 
    2908, 
    2909, 
    2910, 
    2911, 
    2912, 
    2913, 
    2914, 
    2915, 
    2916, 
    2917, 
    2918, 
    2919, 
    2920, 
    2921, 
    2922, 
    2923, 
    2924, 
    2925, 
    2926, 
    2927, 
    2928, 
    2929, 
    2930, 
    2931, 
    2932, 
    2933, 
    2934, 
    2935, 
    2936, 
    2937, 
    2938, 
    2939, 
    2940, 
    2941, 
    2942, 
    2943, 
    2944, 
    2945, 
    2946, 
    2947, 
    2948, 
    2949, 
    2950, 
    2951, 
    2952, 
    2953, 
    2954, 
    2955, 
    2956, 
    2957, 
    2958, 
    2959, 
    2960, 
    2961, 
    2962, 
    2963, 
    2964, 
    2965, 
    2966, 
    2967, 
    2968, 
    2969, 
    2970, 
    2971, 
    2972, 
    2973, 
    2974, 
    2975, 
    2976, 
    2977, 
    2978, 
    2979, 
    2980, 
    2981, 
    2982, 
    2983, 
    2984, 
    2985, 
    2986, 
    2987, 
    2988, 
    2989, 
    2990, 
    2991, 
    2992, 
    2993, 
    2994, 
    2995, 
    2996, 
    2997, 
    2998, 
    2999, 
    3000, 
    3001, 
    3002, 
    3003, 
    3004, 
    3005, 
    3006, 
    3007, 
    3008, 
    3009, 
    3010, 
    3011, 
    3012, 
    3013, 
    3014, 
    3015, 
    3016, 
    3017, 
    3018, 
    3019, 
    3020, 
    3021, 
    3022, 
    3023, 
    3024, 
    3025, 
    3026, 
    3027, 
    3028, 
    3029, 
    3030, 
    3031, 
    3032, 
    3033, 
    3034, 
    3035, 
    3036, 
    3037, 
    3038, 
    3039, 
    3040, 
    3041, 
    3042, 
    3043, 
    3044, 
    3045, 
    3046, 
    3047, 
    3048, 
    3049, 
    3050, 
    3051, 
    3052, 
    3053, 
    3054, 
    3055, 
    3056, 
    3057, 
    3058, 
    3059, 
    3060, 
    3061, 
    3062, 
    3063, 
    3064, 
    3065, 
    3066, 
    3067, 
    3068, 
    3069, 
    3070, 
    3071, 
    3072, 
    3073, 
    3074, 
    3075, 
    3076, 
    3077, 
    3078, 
    3079, 
    3080, 
    3081, 
    3082, 
    3083, 
    3084, 
    3085, 
    3086, 
    3087, 
    3088, 
    3089, 
    3090, 
    3091, 
    3092, 
    3093, 
    3094, 
    3095, 
    3096, 
    3097, 
    3098, 
    3099, 
    3100, 
    3101, 
    3102, 
    3103, 
    3104, 
    3105, 
    3106, 
    3107, 
    3108, 
    3109, 
    3110, 
    3111, 
    3112, 
    3113, 
    3114, 
    3115, 
    3116, 
    3117, 
    3118, 
    3119, 
    3120, 
    3121, 
    3122, 
    3123, 
    3124, 
    3125, 
    3126, 
    3127, 
    3128, 
    3129, 
    3130, 
    3131, 
    3132, 
    3133, 
    3134, 
    3135, 
    3136, 
    3137, 
    3138, 
    3139, 
    3140, 
    3141, 
    3142, 
    3143, 
    3144, 
    3145, 
    3146, 
    3147, 
    3148, 
    3149, 
    3150, 
    3151, 
    3152, 
    3153, 
    3154, 
    3155, 
    3156, 
    3157, 
    3158, 
    3159, 
    3160, 
    3161, 
    3162, 
    3163, 
    3164, 
    3165, 
    3166, 
    3167, 
    3168, 
    3169, 
    3170, 
    3171, 
    3172, 
    3173, 
    3174, 
    3175, 
    3176, 
    3177, 
    3178, 
    3179, 
    3180, 
    3181, 
    3182, 
    3183, 
    3184, 
    3185, 
    3186, 
    3187, 
    3188, 
    3189, 
    3190, 
    3191, 
    3192, 
    3193, 
    3194, 
    3195, 
    3196, 
    3197, 
    3198, 
    3199, 
    3200, 
    3201, 
    3202, 
    3203, 
    3204, 
    3205, 
    3206, 
    3207, 
    3208, 
    3209, 
    3210, 
    3211, 
    3212, 
    3213, 
    3214, 
    3215, 
    3216, 
    3217, 
    3218, 
    3219, 
    3220, 
    3221, 
    3222, 
    3223, 
    3224, 
    3225, 
    3226, 
    3227, 
    3228, 
    3229, 
    3230, 
    3231, 
    3232, 
    3233, 
    3234, 
    3235, 
    3236, 
    3237, 
    3238, 
    3239, 
    3240, 
    3241, 
    3242, 
    3243, 
    3244, 
    3245, 
    3246, 
    3247, 
    3248, 
    3249, 
    3250, 
    3251, 
    3252, 
    3253, 
    3254, 
    3255, 
    3256, 
    3257, 
    3258, 
    3259, 
    3260, 
    3261, 
    3262, 
    3263, 
    3264, 
    3265, 
    3266, 
    3267, 
    3268, 
    3269, 
    3270, 
    3271, 
    3272, 
    3273, 
    3274, 
    3275, 
    3276, 
    3277, 
    3278, 
    3279, 
    3280, 
    3281, 
    3282, 
    3283, 
    3284, 
    3285, 
    3286, 
    3287, 
    3288, 
    3289, 
    3290, 
    3291, 
    3292, 
    3293, 
    3294, 
    3295, 
    3296, 
    3297, 
    3298, 
    3299, 
    3300, 
    3301, 
    3302, 
    3303, 
    3304, 
    3305, 
    3306, 
    3307, 
    3308, 
    3309, 
    3310, 
    3311, 
    3312, 
    3313, 
    3314, 
    3315, 
    3316, 
    3317, 
    3318, 
    3319, 
    3320, 
    3321, 
    3322, 
    3323, 
    3324, 
    3325, 
    3326, 
    3327, 
    3328, 
    3329, 
    3330, 
    3331, 
    3332, 
    3333, 
    3334, 
    3335, 
    3336, 
    3337, 
    3338, 
    3339, 
    3340, 
    3341, 
    3342, 
    3343, 
    3344, 
    3345, 
    3346, 
    3347, 
    3348, 
    3349, 
    3350, 
    3351, 
    3352, 
    3353, 
    3354, 
    3355, 
    3356, 
    3357, 
    3358, 
    3359, 
    3360, 
    3361, 
    3362, 
    3363, 
    3364, 
    3365, 
    3366, 
    3367, 
    3368, 
    3369, 
    3370, 
    3371, 
    3372, 
    3373, 
    3374, 
    3375, 
    3376, 
    3377, 
    3378, 
    3379, 
    3380, 
    3381, 
    3382, 
    3383, 
    3384, 
    3385, 
    3386, 
    3387, 
    3388, 
    3389, 
    3390, 
    3391, 
    3392, 
    3393, 
    3394, 
    3395, 
    3396, 
    3397, 
    3398, 
    3399, 
    3400, 
    3401, 
    3402, 
    3403, 
    3404, 
    3405, 
    3406, 
    3407, 
    3408, 
    3409, 
    3410, 
    3411, 
    3412, 
    3413, 
    3414, 
    3415, 
    3416, 
    3417, 
    3418, 
    3419, 
    3420, 
    3421, 
    3422, 
    3423, 
    3424, 
    3425, 
    3426, 
    3427, 
    3428, 
    3429, 
    3430, 
    3431, 
    3432, 
    3433, 
    3434, 
    3435, 
    3436, 
    3437, 
    3438, 
    3439, 
    3440, 
    3441, 
    3442, 
    3443, 
    3444, 
    3445, 
    3446, 
    3447, 
    3448, 
    3449, 
    3450, 
    3451, 
    3452, 
    3453, 
    3454, 
    3455, 
    3456, 
    3457, 
    3458, 
    3459, 
    3460, 
    3461, 
    3462, 
    3463, 
    3464, 
    3465, 
    3466, 
    3467, 
    3468, 
    3469, 
    3470, 
    3471, 
    3472, 
    3473, 
    3474, 
    3475, 
    3476, 
    3477, 
    3478, 
    3479, 
    3480, 
    3481, 
    3482, 
    3483, 
    3484, 
    3485, 
    3486, 
    3487, 
    3488, 
    3489, 
    3490, 
    3491, 
    3492, 
    3493, 
    3494, 
    3495, 
    3496, 
    3497, 
    3498, 
    3499, 
    3500, 
    3501, 
    3502, 
    3503, 
    3504, 
    3505, 
    3506, 
    3507, 
    3508, 
    3509, 
    3510, 
    3511, 
    3512, 
    3513, 
    3514, 
    3515, 
    3516, 
    3517, 
    3518, 
    3519, 
    3520, 
    3521, 
    3522, 
    3523, 
    3524, 
    3525, 
    3526, 
    3527, 
    3528, 
    3529, 
    3530, 
    3531, 
    3532, 
    3533, 
    3534, 
    3535, 
    3536, 
    3537, 
    3538, 
    3539, 
    3540, 
    3541, 
    3542, 
    3543, 
    3544, 
    3545, 
    3546, 
    3547, 
    3548, 
    3549, 
    3550, 
    3551, 
    3552, 
    3553, 
    3554, 
    3555, 
    3556, 
    3557, 
    3558, 
    3559, 
    3560, 
    3561, 
    3562, 
    3563, 
    3564, 
    3565, 
    3566, 
    3567, 
    3568, 
    3569, 
    3570, 
    3571, 
    3572, 
    3573, 
    3574, 
    3575, 
    3576, 
    3577, 
    3578, 
    3579, 
    3580, 
    3581, 
    3582, 
    3583, 
    3584, 
    3585, 
    3586, 
    3587, 
    3588, 
    3589, 
    3590, 
    3591, 
    3592, 
    3593, 
    3594, 
    3595, 
    3596, 
    3597, 
    3598, 
    3599, 
    3600, 
    3601, 
    3602, 
    3603, 
    3604, 
    3605, 
    3606, 
    3607, 
    3608, 
    3609, 
    3610, 
    3611, 
    3612, 
    3613, 
    3614, 
    3615, 
    3616, 
    3617, 
    3618, 
    3619, 
    3620, 
    3621, 
    3622, 
    3623, 
    3624, 
    3625, 
    3626, 
    3627, 
    3628, 
    3629, 
    3630, 
    3631, 
    3632, 
    3633, 
    3634, 
    3635, 
    3636, 
    3637, 
    3638, 
    3639, 
    3640, 
    3641, 
    3642, 
    3643, 
    3644, 
    3645, 
    3646, 
    3647, 
    3648, 
    3649, 
    3650, 
    3651, 
    3652, 
    3653, 
    3654, 
    3655, 
    3656, 
    3657, 
    3658, 
    3659, 
    3660, 
    3661, 
    3662, 
    3663, 
    3664, 
    3665, 
    3666, 
    3667, 
    3668, 
    3669, 
    3670, 
    3671, 
    3672, 
    3673, 
    3674, 
    3675, 
    3676, 
    3677, 
    3678, 
    3679, 
    3680, 
    3681, 
    3682, 
    3683, 
    3684, 
    3685, 
    3686, 
    3687, 
    3688, 
    3689, 
    3690, 
    3691, 
    3692, 
    3693, 
    3694, 
    3695, 
    3696, 
    3697, 
    3698, 
    3699, 
    3700, 
    3701, 
    3702, 
    3703, 
    3704, 
    3705, 
    3706, 
    3707, 
    3708, 
    3709, 
    3710, 
    3711, 
    3712, 
    3713, 
    3714, 
    3715, 
    3716, 
    3717, 
    3718, 
    3719, 
    3720, 
    3721, 
    3722, 
    3723, 
    3724, 
    3725, 
    3726, 
    3727, 
    3728, 
    3729, 
    3730, 
    3731, 
    3732, 
    3733, 
    3734, 
    3735, 
    3736, 
    3737, 
    3738, 
    3739, 
    3740, 
    3741, 
    3742, 
    3743, 
    3744, 
    3745, 
    3746, 
    3747, 
    3748, 
    3749, 
    3750, 
    3751, 
    3752, 
    3753, 
    3754, 
    3755, 
    3756, 
    3757, 
    3758, 
    3759, 
    3760, 
    3761, 
    3762, 
    3763, 
    3764, 
    3765, 
    3766, 
    3767, 
    3768, 
    3769, 
    3770, 
    3771, 
    3772, 
    3773, 
    3774, 
    3775, 
    3776, 
    3777, 
    3778, 
    3779, 
    3780, 
    3781, 
    3782, 
    3783, 
    3784, 
    3785, 
    3786, 
    3787, 
    3788, 
    3789, 
    3790, 
    3791, 
    3792, 
    3793, 
    3794, 
    3795, 
    3796, 
    3797, 
    3798, 
    3799, 
    3800, 
    3801, 
    3802, 
    3803, 
    3804, 
    3805, 
    3806, 
    3807, 
    3808, 
    3809, 
    3810, 
    3811, 
    3812, 
    3813, 
    3814, 
    3815, 
    3816, 
    3817, 
    3818, 
    3819, 
    3820, 
    3821, 
    3822, 
    3823, 
    3824, 
    3825, 
    3826, 
    3827, 
    3828, 
    3829, 
    3830, 
    3831, 
    3832, 
    3833, 
    3834, 
    3835, 
    3836, 
    3837, 
    3838, 
    3839, 
    3840, 
    3841, 
    3842, 
    3843, 
    3844, 
    3845, 
    3846, 
    3847, 
    3848, 
    3849, 
    3850, 
    3851, 
    3852, 
    3853, 
    3854, 
    3855, 
    3856, 
    3857, 
    3858, 
    3859, 
    3860, 
    3861, 
    3862, 
    3863, 
    3864, 
    3865, 
    3866, 
    3867, 
    3868, 
    3869, 
    3870, 
    3871, 
    3872, 
    3873, 
    3874, 
    3875, 
    3876, 
    3877, 
    3878, 
    3879, 
    3880, 
    3881, 
    3882, 
    3883, 
    3884, 
    3885, 
    3886, 
    3887, 
    3888, 
    3889, 
    3890, 
    3891, 
    3892, 
    3893, 
    3894, 
    3895, 
    3896, 
    3897, 
    3898, 
    3899, 
    3900, 
    3901, 
    3902, 
    3903, 
    3904, 
    3905, 
    3906, 
    3907, 
    3908, 
    3909, 
    3910, 
    3911, 
    3912, 
    3913, 
    3914, 
    3915, 
    3916, 
    3917, 
    3918, 
    3919, 
    3920, 
    3921, 
    3922, 
    3923, 
    3924, 
    3925, 
    3926, 
    3927, 
    3928, 
    3929, 
    3930, 
    3931, 
    3932, 
    3933, 
    3934, 
    3935, 
    3936, 
    3937, 
    3938, 
    3939, 
    3940, 
    3941, 
    3942, 
    3943, 
    3944, 
    3945, 
    3946, 
    3947, 
    3948, 
    3949, 
    3950, 
    3951, 
    3952, 
    3953, 
    3954, 
    3955, 
    3956, 
    3957, 
    3958, 
    3959, 
    3960, 
    3961, 
    3962, 
    3963, 
    3964, 
    3965, 
    3966, 
    3967, 
    3968, 
    3969, 
    3970, 
    3971, 
    3972, 
    3973, 
    3974, 
    3975, 
    3976, 
    3977, 
    3978, 
    3979, 
    3980, 
    3981, 
    3982, 
    3983, 
    3984, 
    3985, 
    3986, 
    3987, 
    3988, 
    3989, 
    3990, 
    3991, 
    3992, 
    3993, 
    3994, 
    3995, 
    3996, 
    3997, 
    3998, 
    3999, 
    4000, 
    4001, 
    4002, 
    4003, 
    4004, 
    4005, 
    4006, 
    4007, 
    4008, 
    4009, 
    4010, 
    4011, 
    4012, 
    4013, 
    4014, 
    4015, 
    4016, 
    4017, 
    4018, 
    4019, 
    4020, 
    4021, 
    4022, 
    4023, 
    4024, 
    4025, 
    4026, 
    4027, 
    4028, 
    4029, 
    4030, 
    4031, 
    4032, 
    4033, 
    4034, 
    4035, 
    4036, 
    4037, 
    4038, 
    4039, 
    4040, 
    4041, 
    4042, 
    4043, 
    4044, 
    4045, 
    4046, 
    4047, 
    4048, 
    4049, 
    4050, 
    4051, 
    4052, 
    4053, 
    4054, 
    4055, 
    4056, 
    4057, 
    4058, 
    4059, 
    4060, 
    4061, 
    4062, 
    4063, 
    4064, 
    4065, 
    4066, 
    4067, 
    4068, 
    4069, 
    4070, 
    4071, 
    4072, 
    4073, 
    4074, 
    4075, 
    4076, 
    4077, 
    4078, 
    4079, 
    4080, 
    4081, 
    4082, 
    4083, 
    4084, 
    4085, 
    4086, 
    4087, 
    4088, 
    4089, 
    4090, 
    4091, 
    4092, 
    4093, 
    4094, 
    4095, 
    4096, 
    4097, 
    4098, 
    4099, 
    4100, 
    4101, 
    4102, 
    4103, 
    4104, 
    4105, 
    4106, 
    4107, 
    4108, 
    4109, 
    4110, 
    4111, 
    4112, 
    4113, 
    4114, 
    4115, 
    4116, 
    4117, 
    4118, 
    4119, 
    4120, 
    4121, 
    4122, 
    4123, 
    4124, 
    4125, 
    4126, 
    4127, 
    4128, 
    4129, 
    4130, 
    4131, 
    4132, 
    4133, 
    4134, 
    4135, 
    4136, 
    4137, 
    4138, 
    4139, 
    4140, 
    4141, 
    4142, 
    4143, 
    4144, 
    4145, 
    4146, 
    4147, 
    4148, 
    4149, 
    4150, 
    4151, 
    4152, 
    4153, 
    4154, 
    4155, 
    4156, 
    4157, 
    4158, 
    4159, 
    4160, 
    4161, 
    4162, 
    4163, 
    4164, 
    4165, 
    4166, 
    4167, 
    4168, 
    4169, 
    4170, 
    4171, 
    4172, 
    4173, 
    4174, 
    4175, 
    4176, 
    4177, 
    4178, 
    4179, 
    4180, 
    4181, 
    4182, 
    4183, 
    4184, 
    4185, 
    4186, 
    4187, 
    4188, 
    4189, 
    4190, 
    4191, 
    4192, 
    4193, 
    4194, 
    4195, 
    4196, 
    4197, 
    4198, 
    4199, 
    4200, 
    4201, 
    4202, 
    4203, 
    4204, 
    4205, 
    4206, 
    4207, 
    4208, 
    4209, 
    4210, 
    4211, 
    4212, 
    4213, 
    4214, 
    4215, 
    4216, 
    4217, 
    4218, 
    4219, 
    4220, 
    4221, 
    4222, 
    4223, 
    4224, 
    4225, 
    4226, 
    4227, 
    4228, 
    4229, 
    4230, 
    4231, 
    4232, 
    4233, 
    4234, 
    4235, 
    4236, 
    4237, 
    4238, 
    4239, 
    4240, 
    4241, 
    4242, 
    4243, 
    4244, 
    4245, 
    4246, 
    4247, 
    4248, 
    4249, 
    4250, 
    4251, 
    4252, 
    4253, 
    4254, 
    4255, 
    4256, 
    4257, 
    4258, 
    4259, 
    4260, 
    4261, 
    4262, 
    4263, 
    4264, 
    4265, 
    4266, 
    4267, 
    4268, 
    4269, 
    4270, 
    4271, 
    4272, 
    4273, 
    4274, 
    4275, 
    4276, 
    4277, 
    4278, 
    4279, 
    4280, 
    4281, 
    4282, 
    4283, 
    4284, 
    4285, 
    4286, 
    4287, 
    4288, 
    4289, 
    4290, 
    4291, 
    4292, 
    4293, 
    4294, 
    4295, 
    4296, 
    4297, 
    4298, 
    4299, 
    4300, 
    4301, 
    4302, 
    4303, 
    4304, 
    4305, 
    4306, 
    4307, 
    4308, 
    4309, 
    4310, 
    4311, 
    4312, 
    4313, 
    4314, 
    4315, 
    4316, 
    4317, 
    4318, 
    4319, 
    4320, 
    4321, 
    4322, 
    4323, 
    4324, 
    4325, 
    4326, 
    4327, 
    4328, 
    4329, 
    4330, 
    4331, 
    4332, 
    4333, 
    4334, 
    4335, 
    4336, 
    4337, 
    4338, 
    4339, 
    4340, 
    4341, 
    4342, 
    4343, 
    4344, 
    4345, 
    4346, 
    4347, 
    4348, 
    4349, 
    4350, 
    4351, 
    4352, 
    4353, 
    4354, 
    4355, 
    4356, 
    4357, 
    4358, 
    4359, 
    4360, 
    4361, 
    4362, 
    4363, 
    4364, 
    4365, 
    4366, 
    4367, 
    4368, 
    4369, 
    4370, 
    4371, 
    4372, 
    4373, 
    4374, 
    4375, 
    4376, 
    4377, 
    4378, 
    4379, 
    4380, 
    4381, 
    4382, 
    4383, 
    4384, 
    4385, 
    4386, 
    4387, 
    4388, 
    4389, 
    4390, 
    4391, 
    4392, 
    4393, 
    4394, 
    4395, 
    4396, 
    4397, 
    4398, 
    4399, 
    4400, 
    4401, 
    4402, 
    4403, 
    4404, 
    4405, 
    4406, 
    4407, 
    4408, 
    4409, 
    4410, 
    4411, 
    4412, 
    4413, 
    4414, 
    4415, 
    4416, 
    4417, 
    4418, 
    4419, 
    4420, 
    4421, 
    4422, 
    4423, 
    4424, 
    4425, 
    4426, 
    4427, 
    4428, 
    4429, 
    4430, 
    4431, 
    4432, 
    4433, 
    4434, 
    4435, 
    4436, 
    4437, 
    4438, 
    4439, 
    4440, 
    4441, 
    4442, 
    4443, 
    4444, 
    4445, 
    4446, 
    4447, 
    4448, 
    4449, 
    4450, 
    4451, 
    4452, 
    4453, 
    4454, 
    4455, 
    4456, 
    4457, 
    4458, 
    4459, 
    4460, 
    4461, 
    4462, 
    4463, 
    4464, 
    4465, 
    4466, 
    4467, 
    4468, 
    4469, 
    4470, 
    4471, 
    4472, 
    4473, 
    4474, 
    4475, 
    4476, 
    4477, 
    4478, 
    4479, 
    4480, 
    4481, 
    4482, 
    4483, 
    4484, 
    4485, 
    4486, 
    4487, 
    4488, 
    4489, 
    4490, 
    4491, 
    4492, 
    4493, 
    4494, 
    4495, 
    4496, 
    4497, 
    4498, 
    4499, 
    4500, 
    4501, 
    4502, 
    4503, 
    4504, 
    4505, 
    4506, 
    4507, 
    4508, 
    4509, 
    4510, 
    4511, 
    4512, 
    4513, 
    4514, 
    4515, 
    4516, 
    4517, 
    4518, 
    4519, 
    4520, 
    4521, 
    4522, 
    4523, 
    4524, 
    4525, 
    4526, 
    4527, 
    4528, 
    4529, 
    4530, 
    4531, 
    4532, 
    4533, 
    4534, 
    4535, 
    4536, 
    4537, 
    4538, 
    4539, 
    4540, 
    4541, 
    4542, 
    4543, 
    4544, 
    4545, 
    4546, 
    4547, 
    4548, 
    4549, 
    4550, 
    4551, 
    4552, 
    4553, 
    4554, 
    4555, 
    4556, 
    4557, 
    4558, 
    4559, 
    4560, 
    4561, 
    4562, 
    4563, 
    4564, 
    4565, 
    4566, 
    4567, 
    4568, 
    4569, 
    4570, 
    4571, 
    4572, 
    4573, 
    4574, 
    4575, 
    4576, 
    4577, 
    4578, 
    4579, 
    4580, 
    4581, 
    4582, 
    4583, 
    4584, 
    4585, 
    4586, 
    4587, 
    4588, 
    4589, 
    4590, 
    4591, 
    4592, 
    4593, 
    4594, 
    4595, 
    4596, 
    4597, 
    4598, 
    4599, 
    4600, 
    4601, 
    4602, 
    4603, 
    4604, 
    4605, 
    4606, 
    4607, 
    4608, 
    4609, 
    4610, 
    4611, 
    4612, 
    4613, 
    4614, 
    4615, 
    4616, 
    4617, 
    4618, 
    4619, 
    4620, 
    4621, 
    4622, 
    4623, 
    4624, 
    4625, 
    4626, 
    4627, 
    4628, 
    4629, 
    4630, 
    4631, 
    4632, 
    4633, 
    4634, 
    4635, 
    4636, 
    4637, 
    4638, 
    4639, 
    4640, 
    4641, 
    4642, 
    4643, 
    4644, 
    4645, 
    4646, 
    4647, 
    4648, 
    4649, 
    4650, 
    4651, 
    4652, 
    4653, 
    4654, 
    4655, 
    4656, 
    4657, 
    4658, 
    4659, 
    4660, 
    4661, 
    4662, 
    4663, 
    4664, 
    4665, 
    4666, 
    4667, 
    4668, 
    4669, 
    4670, 
    4671, 
    4672, 
    4673, 
    4674, 
    4675, 
    4676, 
    4677, 
    4678, 
    4679, 
    4680, 
    4681, 
    4682, 
    4683, 
    4684, 
    4685, 
    4686, 
    4687, 
    4688, 
    4689, 
    4690, 
    4691, 
    4692, 
    4693, 
    4694, 
    4695, 
    4696, 
    4697, 
    4698, 
    4699, 
    4700, 
    4701, 
    4702, 
    4703, 
    4704, 
    4705, 
    4706, 
    4707, 
    4708, 
    4709, 
    4710, 
    4711, 
    4712, 
    4713, 
    4714, 
    4715, 
    4716, 
    4717, 
    4718, 
    4719, 
    4720, 
    4721, 
    4722, 
    4723, 
    4724, 
    4725, 
    4726, 
    4727, 
    4728, 
    4729, 
    4730, 
    4731, 
    4732, 
    4733, 
    4734, 
    4735, 
    4736, 
    4737, 
    4738, 
    4739, 
    4740, 
    4741, 
    4742, 
    4743, 
    4744, 
    4745, 
    4746, 
    4747, 
    4748, 
    4749, 
    4750, 
    4751, 
    4752, 
    4753, 
    4754, 
    4755, 
    4756, 
    4757, 
    4758, 
    4759, 
    4760, 
    4761, 
    4762, 
    4763, 
    4764, 
    4765, 
    4766, 
    4767, 
    4768, 
    4769, 
    4770, 
    4771, 
    4772, 
    4773, 
    4774, 
    4775, 
    4776, 
    4777, 
    4778, 
    4779, 
    4780, 
    4781, 
    4782, 
    4783, 
    4784, 
    4785, 
    4786, 
    4787, 
    4788, 
    4789, 
    4790, 
    4791, 
    4792, 
    4793, 
    4794, 
    4795, 
    4796, 
    4797, 
    4798, 
    4799, 
    4800, 
    4801, 
    4802, 
    4803, 
    4804, 
    4805, 
    4806, 
    4807, 
    4808, 
    4809, 
    4810, 
    4811, 
    4812, 
    4813, 
    4814, 
    4815, 
    4816, 
    4817, 
    4818, 
    4819, 
    4820, 
    4821, 
    4822, 
    4823, 
    4824, 
    4825, 
    4826, 
    4827, 
    4828, 
    4829, 
    4830, 
    4831, 
    4832, 
    4833, 
    4834, 
    4835, 
    4836, 
    4837, 
    4838, 
    4839, 
    4840, 
    4841, 
    4842, 
    4843, 
    4844, 
    4845, 
    4846, 
    4847, 
    4848, 
    4849, 
    4850, 
    4851, 
    4852, 
    4853, 
    4854, 
    4855, 
    4856, 
    4857, 
    4858, 
    4859, 
    4860, 
    4861, 
    4862, 
    4863, 
    4864, 
    4865, 
    4866, 
    4867, 
    4868, 
    4869, 
    4870, 
    4871, 
    4872, 
    4873, 
    4874, 
    4875, 
    4876, 
    4877, 
    4878, 
    4879, 
    4880, 
    4881, 
    4882, 
    4883, 
    4884, 
    4885, 
    4886, 
    4887, 
    4888, 
    4889, 
    4890, 
    4891, 
    4892, 
    4893, 
    4894, 
    4895, 
    4896, 
    4897, 
    4898, 
    4899, 
    4900, 
    4901, 
    4902, 
    4903, 
    4904, 
    4905, 
    4906, 
    4907, 
    4908, 
    4909, 
    4910, 
    4911, 
    4912, 
    4913, 
    4914, 
    4915, 
    4916, 
    4917, 
    4918, 
    4919, 
    4920, 
    4921, 
    4922, 
    4923, 
    4924, 
    4925, 
    4926, 
    4927, 
    4928, 
    4929, 
    4930, 
    4931, 
    4932, 
    4933, 
    4934, 
    4935, 
    4936, 
    4937, 
    4938, 
    4939, 
    4940, 
    4941, 
    4942, 
    4943, 
    4944, 
    4945, 
    4946, 
    4947, 
    4948, 
    4949, 
    4950, 
    4951, 
    4952, 
    4953, 
    4954, 
    4955, 
    4956, 
    4957, 
    4958, 
    4959, 
    4960, 
    4961, 
    4962, 
    4963, 
    4964, 
    4965, 
    4966, 
    4967, 
    4968, 
    4969, 
    4970, 
    4971, 
    4972, 
    4973, 
    4974, 
    4975, 
    4976, 
    4977, 
    4978, 
    4979, 
    4980, 
    4981, 
    4982, 
    4983, 
    4984, 
    4985, 
    4986, 
    4987, 
    4988, 
    4989, 
    4990, 
    4991, 
    4992, 
    4993, 
    4994, 
    4995, 
    4996, 
    4997, 
    4998, 
    4999, 
    5000, 
    5001, 
    5002, 
    5003, 
    5004, 
    5005, 
    5006, 
    5007, 
    5008, 
    5009, 
    5010, 
    5011, 
    5012, 
    5013, 
    5014, 
    5015, 
    5016, 
    5017, 
    5018, 
    5019, 
    5020, 
    5021, 
    5022, 
    5023, 
    5024, 
    5025, 
    5026, 
    5027, 
    5028, 
    5029, 
    5030, 
    5031, 
    5032, 
    5033, 
    5034, 
    5035, 
    5036, 
    5037, 
    5038, 
    5039, 
    5040, 
    5041, 
    5042, 
    5043, 
    5044, 
    5045, 
    5046, 
    5047, 
    5048, 
    5049, 
    5050, 
    5051, 
    5052, 
    5053, 
    5054, 
    5055, 
    5056, 
    5057, 
    5058, 
    5059, 
    5060, 
    5061, 
    5062, 
    5063, 
    5064, 
    5065, 
    5066, 
    5067, 
    5068, 
    5069, 
    5070, 
    5071, 
    5072, 
    5073, 
    5074, 
    5075, 
    5076, 
    5077, 
    5078, 
    5079, 
    5080, 
    5081, 
    5082, 
    5083, 
    5084, 
    5085, 
    5086, 
    5087, 
    5088, 
    5089, 
    5090, 
    5091, 
    5092, 
    5093, 
    5094, 
    5095, 
    5096, 
    5097, 
    5098, 
    5099, 
    5100, 
    5101, 
    5102, 
    5103, 
    5104, 
    5105, 
    5106, 
    5107, 
    5108, 
    5109, 
    5110, 
    5111, 
    5112, 
    5113, 
    5114, 
    5115, 
    5116, 
    5117, 
    5118, 
    5119, 
    5120, 
    5121, 
    5122, 
    5123, 
    5124, 
    5125, 
    5126, 
    5127, 
    5128, 
    5129, 
    5130, 
    5131, 
    5132, 
    5133, 
    5134, 
    5135, 
    5136, 
    5137, 
    5138, 
    5139, 
    5140, 
    5141, 
    5142, 
    5143, 
    5144, 
    5145, 
    5146, 
    5147, 
    5148, 
    5149, 
    5150, 
    5151, 
    5152, 
    5153, 
    5154, 
    5155, 
    5156, 
    5157, 
    5158, 
    5159, 
    5160, 
    5161, 
    5162, 
    5163, 
    5164, 
    5165, 
    5166, 
    5167, 
    5168, 
    5169, 
    5170, 
    5171, 
    5172, 
    5173, 
    5174, 
    5175, 
    5176, 
    5177, 
    5178, 
    5179, 
    5180, 
    5181, 
    5182, 
    5183, 
    5184, 
    5185, 
    5186, 
    5187, 
    5188, 
    5189, 
    5190, 
    5191, 
    5192, 
    5193, 
    5194, 
    5195, 
    5196, 
    5197, 
    5198, 
    5199, 
    5200, 
    5201, 
    5202, 
    5203, 
    5204, 
    5205, 
    5206, 
    5207, 
    5208, 
    5209, 
    5210, 
    5211, 
    5212, 
    5213, 
    5214, 
    5215, 
    5216, 
    5217, 
    5218, 
    5219, 
    5220, 
    5221, 
    5222, 
    5223, 
    5224, 
    5225, 
    5226, 
    5227, 
    5228, 
    5229, 
    5230, 
    5231, 
    5232, 
    5233, 
    5234, 
    5235, 
    5236, 
    5237, 
    5238, 
    5239, 
    5240, 
    5241, 
    5242, 
    5243, 
    5244, 
    5245, 
    5246, 
    5247, 
    5248, 
    5249, 
    5250, 
    5251, 
    5252, 
    5253, 
    5254, 
    5255, 
    5256, 
    5257, 
    5258, 
    5259, 
    5260, 
    5261, 
    5262, 
    5263, 
    5264, 
    5265, 
    5266, 
    5267, 
    5268, 
    5269, 
    5270, 
    5271, 
    5272, 
    5273, 
    5274, 
    5275, 
    5276, 
    5277, 
    5278, 
    5279, 
    5280, 
    5281, 
    5282, 
    5283, 
    5284, 
    5285, 
    5286, 
    5287, 
    5288, 
    5289, 
    5290, 
    5291, 
    5292, 
    5293, 
    5294, 
    5295, 
    5296, 
    5297, 
    5298, 
    5299, 
    5300, 
    5301, 
    5302, 
    5303, 
    5304, 
    5305, 
    5306, 
    5307, 
    5308, 
    5309, 
    5310, 
    5311, 
    5312, 
    5313, 
    5314, 
    5315, 
    5316, 
    5317, 
    5318, 
    5319, 
    5320, 
    5321, 
    5322, 
    5323, 
    5324, 
    5325, 
    5326, 
    5327, 
    5328, 
    5329, 
    5330, 
    5331, 
    5332, 
    5333, 
    5334, 
    5335, 
    5336, 
    5337, 
    5338, 
    5339, 
    5340, 
    5341, 
    5342, 
    5343, 
    5344, 
    5345, 
    5346, 
    5347, 
    5348, 
    5349, 
    5350, 
    5351, 
    5352, 
    5353, 
    5354, 
    5355, 
    5356, 
    5357, 
    5358, 
    5359, 
    5360, 
    5361, 
    5362, 
    5363, 
    5364, 
    5365, 
    5366, 
    5367, 
    5368, 
    5369, 
    5370, 
    5371, 
    5372, 
    5373, 
    5374, 
    5375, 
    5376, 
    5377, 
    5378, 
    5379, 
    5380, 
    5381, 
    5382, 
    5383, 
    5384, 
    5385, 
    5386, 
    5387, 
    5388, 
    5389, 
    5390, 
    5391, 
    5392, 
    5393, 
    5394, 
    5395, 
    5396, 
    5397, 
    5398, 
    5399, 
    5400, 
    5401, 
    5402, 
    5403, 
    5404, 
    5405, 
    5406, 
    5407, 
    5408, 
    5409, 
    5410, 
    5411, 
    5412, 
    5413, 
    5414, 
    5415, 
    5416, 
    5417, 
    5418, 
    5419, 
    5420, 
    5421, 
    5422, 
    5423, 
    5424, 
    5425, 
    5426, 
    5427, 
    5428, 
    5429, 
    5430, 
    5431, 
    5432, 
    5433, 
    5434, 
    5435, 
    5436, 
    5437, 
    5438, 
    5439, 
    5440, 
    5441, 
    5442, 
    5443, 
    5444, 
    5445, 
    5446, 
    5447, 
    5448, 
    5449, 
    5450, 
    5451, 
    5452, 
    5453, 
    5454, 
    5455, 
    5456, 
    5457, 
    5458, 
    5459, 
    5460, 
    5461, 
    5462, 
    5463, 
    5464, 
    5465, 
    5466, 
    5467, 
    5468, 
    5469, 
    5470, 
    5471, 
    5472, 
    5473, 
    5474, 
    5475, 
    5476, 
    5477, 
    5478, 
    5479, 
    5480, 
    5481, 
    5482, 
    5483, 
    5484, 
    5485, 
    5486, 
    5487, 
    5488, 
    5489, 
    5490, 
    5491, 
    5492, 
    5493, 
    5494, 
    5495, 
    5496, 
    5497, 
    5498, 
    5499, 
    5500, 
    5501, 
    5502, 
    5503, 
    5504, 
    5505, 
    5506, 
    5507, 
    5508, 
    5509, 
    5510, 
    5511, 
    5512, 
    5513, 
    5514, 
    5515, 
    5516, 
    5517, 
    5518, 
    5519, 
    5520, 
    5521, 
    5522, 
    5523, 
    5524, 
    5525, 
    5526, 
    5527, 
    5528, 
    5529, 
    5530, 
    5531, 
    5532, 
    5533, 
    5534, 
    5535, 
    5536, 
    5537, 
    5538, 
    5539, 
    5540, 
    5541, 
    5542, 
    5543, 
    5544, 
    5545, 
    5546, 
    5547, 
    5548, 
    5549, 
    5550, 
    5551, 
    5552, 
    5553, 
    5554, 
    5555, 
    5556, 
    5557, 
    5558, 
    5559, 
    5560, 
    5561, 
    5562, 
    5563, 
    5564, 
    5565, 
    5566, 
    5567, 
    5568, 
    5569, 
    5570, 
    5571, 
    5572, 
    5573, 
    5574, 
    5575, 
    5576, 
    5577, 
    5578, 
    5579, 
    5580, 
    5581, 
    5582, 
    5583, 
    5584, 
    5585, 
    5586, 
    5587, 
    5588, 
    5589, 
    5590, 
    5591, 
    5592, 
    5593, 
    5594, 
    5595, 
    5596, 
    5597, 
    5598, 
    5599, 
    5600, 
    5601, 
    5602, 
    5603, 
    5604, 
    5605, 
    5606, 
    5607, 
    5608, 
    5609, 
    5610, 
    5611, 
    5612, 
    5613, 
    5614, 
    5615, 
    5616, 
    5617, 
    5618, 
    5619, 
    5620, 
    5621, 
    5622, 
    5623, 
    5624, 
    5625, 
    5626, 
    5627, 
    5628, 
    5629, 
    5630, 
    5631, 
    5632, 
    5633, 
    5634, 
    5635, 
    5636, 
    5637, 
    5638, 
    5639, 
    5640, 
    5641, 
    5642, 
    5643, 
    5644, 
    5645, 
    5646, 
    5647, 
    5648, 
    5649, 
    5650, 
    5651, 
    5652, 
    5653, 
    5654, 
    5655, 
    5656, 
    5657, 
    5658, 
    5659, 
    5660, 
    5661, 
    5662, 
    5663, 
    5664, 
    5665, 
    5666, 
    5667, 
    5668, 
    5669, 
    5670, 
    5671, 
    5672, 
    5673, 
    5674, 
    5675, 
    5676, 
    5677, 
    5678, 
    5679, 
    5680, 
    5681, 
    5682, 
    5683, 
    5684, 
    5685, 
    5686, 
    5687, 
    5688, 
    5689, 
    5690, 
    5691, 
    5692, 
    5693, 
    5694, 
    5695, 
    5696, 
    5697, 
    5698, 
    5699, 
    5700, 
    5701, 
    5702, 
    5703, 
    5704, 
    5705, 
    5706, 
    5707, 
    5708, 
    5709, 
    5710, 
    5711, 
    5712, 
    5713, 
    5714, 
    5715, 
    5716, 
    5717, 
    5718, 
    5719, 
    5720, 
    5721, 
    5722, 
    5723, 
    5724, 
    5725, 
    5726, 
    5727, 
    5728, 
    5729, 
    5730, 
    5731, 
    5732, 
    5733, 
    5734, 
    5735, 
    5736, 
    5737, 
    5738, 
    5739, 
    5740, 
    5741, 
    5742, 
    5743, 
    5744, 
    5745, 
    5746, 
    5747, 
    5748, 
    5749, 
    5750, 
    5751, 
    5752, 
    5753, 
    5754, 
    5755, 
    5756, 
    5757, 
    5758, 
    5759, 
    5760, 
    5761, 
    5762, 
    5763, 
    5764, 
    5765, 
    5766, 
    5767, 
    5768, 
    5769, 
    5770, 
    5771, 
    5772, 
    5773, 
    5774, 
    5775, 
    5776, 
    5777, 
    5778, 
    5779, 
    5780, 
    5781, 
    5782, 
    5783, 
    5784, 
    5785, 
    5786, 
    5787, 
    5788, 
    5789, 
    5790, 
    5791, 
    5792, 
    5793, 
    5794, 
    5795, 
    5796, 
    5797, 
    5798, 
    5799, 
    5800, 
    5801, 
    5802, 
    5803, 
    5804, 
    5805, 
    5806, 
    5807, 
    5808, 
    5809, 
    5810, 
    5811, 
    5812, 
    5813, 
    5814, 
    5815, 
    5816, 
    5817, 
    5818, 
    5819, 
    5820, 
    5821, 
    5822, 
    5823, 
    5824, 
    5825, 
    5826, 
    5827, 
    5828, 
    5829, 
    5830, 
    5831, 
    5832, 
    5833, 
    5834, 
    5835, 
    5836, 
    5837, 
    5838, 
    5839, 
    5840, 
    5841, 
    5842, 
    5843, 
    5844, 
    5845, 
    5846, 
    5847, 
    5848, 
    5849, 
    5850, 
    5851, 
    5852, 
    5853, 
    5854, 
    5855, 
    5856, 
    5857, 
    5858, 
    5859, 
    5860, 
    5861, 
    5862, 
    5863, 
    5864, 
    5865, 
    5866, 
    5867, 
    5868, 
    5869, 
    5870, 
    5871, 
    5872, 
    5873, 
    5874, 
    5875, 
    5876, 
    5877, 
    5878, 
    5879, 
    5880, 
    5881, 
    5882, 
    5883, 
    5884, 
    5885, 
    5886, 
    5887, 
    5888, 
    5889, 
    5890, 
    5891, 
    5892, 
    5893, 
    5894, 
    5895, 
    5896, 
    5897, 
    5898, 
    5899, 
    5900, 
    5901, 
    5902, 
    5903, 
    5904, 
    5905, 
    5906, 
    5907, 
    5908, 
    5909, 
    5910, 
    5911, 
    5912, 
    5913, 
    5914, 
    5915, 
    5916, 
    5917, 
    5918, 
    5919, 
    5920, 
    5921, 
    5922, 
    5923, 
    5924, 
    5925, 
    5926, 
    5927, 
    5928, 
    5929, 
    5930, 
    5931, 
    5932, 
    5933, 
    5934, 
    5935, 
    5936, 
    5937, 
    5938, 
    5939, 
    5940, 
    5941, 
    5942, 
    5943, 
    5944, 
    5945, 
    5946, 
    5947, 
    5948, 
    5949, 
    5950, 
    5951, 
    5952, 
    5953, 
    5954, 
    5955, 
    5956, 
    5957, 
    5958, 
    5959, 
    5960, 
    5961, 
    5962, 
    5963, 
    5964, 
    5965, 
    5966, 
    5967, 
    5968, 
    5969, 
    5970, 
    5971, 
    5972, 
    5973, 
    5974, 
    5975, 
    5976, 
    5977, 
    5978, 
    5979, 
    5980, 
    5981, 
    5982, 
    5983, 
    5984, 
    5985, 
    5986, 
    5987, 
    5988, 
    5989, 
    5990, 
    5991, 
    5992, 
    5993, 
    5994, 
    5995, 
    5996, 
    5997, 
    5998, 
    5999, 
    6000, 
    6001, 
    6002, 
    6003, 
    6004, 
    6005, 
    6006, 
    6007, 
    6008, 
    6009, 
    6010, 
    6011, 
    6012, 
    6013, 
    6014, 
    6015, 
    6016, 
    6017, 
    6018, 
    6019, 
    6020, 
    6021, 
    6022, 
    6023, 
    6024, 
    6025, 
    6026, 
    6027, 
    6028, 
    6029, 
    6030, 
    6031, 
    6032, 
    6033, 
    6034, 
    6035, 
    6036, 
    6037, 
    6038, 
    6039, 
    6040, 
    6041, 
    6042, 
    6043, 
    6044, 
    6045, 
    6046, 
    6047, 
    6048, 
    6049, 
    6050, 
    6051, 
    6052, 
    6053, 
    6054, 
    6055, 
    6056, 
    6057, 
    6058, 
    6059, 
    6060, 
    6061, 
    6062, 
    6063, 
    6064, 
    6065, 
    6066, 
    6067, 
    6068, 
    6069, 
    6070, 
    6071, 
    6072, 
    6073, 
    6074, 
    6075, 
    6076, 
    6077, 
    6078, 
    6079, 
    6080, 
    6081, 
    6082, 
    6083, 
    6084, 
    6085, 
    6086, 
    6087, 
    6088, 
    6089, 
    6090, 
    6091, 
    6092, 
    6093, 
    6094, 
    6095, 
    6096, 
    6097, 
    6098, 
    6099, 
    6100, 
    6101, 
    6102, 
    6103, 
    6104, 
    6105, 
    6106, 
    6107, 
    6108, 
    6109, 
    6110, 
    6111, 
    6112, 
    6113, 
    6114, 
    6115, 
    6116, 
    6117, 
    6118, 
    6119, 
    6120, 
    6121, 
    6122, 
    6123, 
    6124, 
    6125, 
    6126, 
    6127, 
    6128, 
    6129, 
    6130, 
    6131, 
    6132, 
    6133, 
    6134, 
    6135, 
    6136, 
    6137, 
    6138, 
    6139, 
    6140, 
    6141, 
    6142, 
    6143, 
    6144, 
    6145, 
    6146, 
    6147, 
    6148, 
    6149, 
    6150, 
    6151, 
    6152, 
    6153, 
    6154, 
    6155, 
    6156, 
    6157, 
    6158, 
    6159, 
    6160, 
    6161, 
    6162, 
    6163, 
    6164, 
    6165, 
    6166, 
    6167, 
    6168, 
    6169, 
    6170, 
    6171, 
    6172, 
    6173, 
    6174, 
    6175, 
    6176, 
    6177, 
    6178, 
    6179, 
    6180, 
    6181, 
    6182, 
    6183, 
    6184, 
    6185, 
    6186, 
    6187, 
    6188, 
    6189, 
    6190, 
    6191, 
    6192, 
    6193, 
    6194, 
    6195, 
    6196, 
    6197, 
    6198, 
    6199, 
    6200, 
    6201, 
    6202, 
    6203, 
    6204, 
    6205, 
    6206, 
    6207, 
    6208, 
    6209, 
    6210, 
    6211, 
    6212, 
    6213, 
    6214, 
    6215, 
    6216, 
    6217, 
    6218, 
    6219, 
    6220, 
    6221, 
    6222, 
    6223, 
    6224, 
    6225, 
    6226, 
    6227, 
    6228, 
    6229, 
    6230, 
    6231, 
    6232, 
    6233, 
    6234, 
    6235, 
    6236, 
    6237, 
    6238, 
    6239, 
    6240, 
    6241, 
    6242, 
    6243, 
    6244, 
    6245, 
    6246, 
    6247, 
    6248, 
    6249, 
    6250, 
    6251, 
    6252, 
    6253, 
    6254, 
    6255, 
    6256, 
    6257, 
    6258, 
    6259, 
    6260, 
    6261, 
    6262, 
    6263, 
    6264, 
    6265, 
    6266, 
    6267, 
    6268, 
    6269, 
    6270, 
    6271, 
    6272, 
    6273, 
    6274, 
    6275, 
    6276, 
    6277, 
    6278, 
    6279, 
    6280, 
    6281, 
    6282, 
    6283, 
    6284, 
    6285, 
    6286, 
    6287, 
    6288, 
    6289, 
    6290, 
    6291, 
    6292, 
    6293, 
    6294, 
    6295, 
    6296, 
    6297, 
    6298, 
    6299, 
    6300, 
    6301, 
    6302, 
    6303, 
    6304, 
    6305, 
    6306, 
    6307, 
    6308, 
    6309, 
    6310, 
    6311, 
    6312, 
    6313, 
    6314, 
    6315, 
    6316, 
    6317, 
    6318, 
    6319, 
    6320, 
    6321, 
    6322, 
    6323, 
    6324, 
    6325, 
    6326, 
    6327, 
    6328, 
    6329, 
    6330, 
    6331, 
    6332, 
    6333, 
    6334, 
    6335, 
    6336, 
    6337, 
    6338, 
    6339, 
    6340, 
    6341, 
    6342, 
    6343, 
    6344, 
    6345, 
    6346, 
    6347, 
    6348, 
    6349, 
    6350, 
    6351, 
    6352, 
    6353, 
    6354, 
    6355, 
    6356, 
    6357, 
    6358, 
    6359, 
    6360, 
    6361, 
    6362, 
    6363, 
    6364, 
    6365, 
    6366, 
    6367, 
    6368, 
    6369, 
    6370, 
    6371, 
    6372, 
    6373, 
    6374, 
    6375, 
    6376, 
    6377, 
    6378, 
    6379, 
    6380, 
    6381, 
    6382, 
    6383, 
    6384, 
    6385, 
    6386, 
    6387, 
    6388, 
    6389, 
    6390, 
    6391, 
    6392, 
    6393, 
    6394, 
    6395, 
    6396, 
    6397, 
    6398, 
    6399, 
    6400, 
    6401, 
    6402, 
    6403, 
    6404, 
    6405, 
    6406, 
    6407, 
    6408, 
    6409, 
    6410, 
    6411, 
    6412, 
    6413, 
    6414, 
    6415, 
    6416, 
    6417, 
    6418, 
    6419, 
    6420, 
    6421, 
    6422, 
    6423, 
    6424, 
    6425, 
    6426, 
    6427, 
    6428, 
    6429, 
    6430, 
    6431, 
    6432, 
    6433, 
    6434, 
    6435, 
    6436, 
    6437, 
    6438, 
    6439, 
    6440, 
    6441, 
    6442, 
    6443, 
    6444, 
    6445, 
    6446, 
    6447, 
    6448, 
    6449, 
    6450, 
    6451, 
    6452, 
    6453, 
    6454, 
    6455, 
    6456, 
    6457, 
    6458, 
    6459, 
    6460, 
    6461, 
    6462, 
    6463, 
    6464, 
    6465, 
    6466, 
    6467, 
    6468, 
    6469, 
    6470, 
    6471, 
    6472, 
    6473, 
    6474, 
    6475, 
    6476, 
    6477, 
    6478, 
    6479, 
    6480, 
    6481, 
    6482, 
    6483, 
    6484, 
    6485, 
    6486, 
    6487, 
    6488, 
    6489, 
    6490, 
    6491, 
    6492, 
    6493, 
    6494, 
    6495, 
    6496, 
    6497, 
    6498, 
    6499, 
    6500, 
    6501, 
    6502, 
    6503, 
    6504, 
    6505, 
    6506, 
    6507, 
    6508, 
    6509, 
    6510, 
    6511, 
    6512, 
    6513, 
    6514, 
    6515, 
    6516, 
    6517, 
    6518, 
    6519, 
    6520, 
    6521, 
    6522, 
    6523, 
    6524, 
    6525, 
    6526, 
    6527, 
    6528, 
    6529, 
    6530, 
    6531, 
    6532, 
    6533, 
    6534, 
    6535, 
    6536, 
    6537, 
    6538, 
    6539, 
    6540, 
    6541, 
    6542, 
    6543, 
    6544, 
    6545, 
    6546, 
    6547, 
    6548, 
    6549, 
    6550, 
    6551, 
    6552, 
    6553, 
    6554, 
    6555, 
    6556, 
    6557, 
    6558, 
    6559, 
    6560, 
    6561, 
    6562, 
    6563, 
    6564, 
    6565, 
    6566, 
    6567, 
    6568, 
    6569, 
    6570, 
    6571, 
    6572, 
    6573, 
    6574, 
    6575, 
    6576, 
    6577, 
    6578, 
    6579, 
    6580, 
    6581, 
    6582, 
    6583, 
    6584, 
    6585, 
    6586, 
    6587, 
    6588, 
    6589, 
    6590, 
    6591, 
    6592, 
    6593, 
    6594, 
    6595, 
    6596, 
    6597, 
    6598, 
    6599, 
    6600, 
    6601, 
    6602, 
    6603, 
    6604, 
    6605, 
    6606, 
    6607, 
    6608, 
    6609, 
    6610, 
    6611, 
    6612, 
    6613, 
    6614, 
    6615, 
    6616, 
    6617, 
    6618, 
    6619, 
    6620, 
    6621, 
    6622, 
    6623, 
    6624, 
    6625, 
    6626, 
    6627, 
    6628, 
    6629, 
    6630, 
    6631, 
    6632, 
    6633, 
    6634, 
    6635, 
    6636, 
    6637, 
    6638, 
    6639, 
    6640, 
    6641, 
    6642, 
    6643, 
    6644, 
    6645, 
    6646, 
    6647, 
    6648, 
    6649, 
    6650, 
    6651, 
    6652, 
    6653, 
    6654, 
    6655, 
    6656, 
    6657, 
    6658, 
    6659, 
    6660, 
    6661, 
    6662, 
    6663, 
    6664, 
    6665, 
    6666, 
    6667, 
    6668, 
    6669, 
    6670, 
    6671, 
    6672, 
    6673, 
    6674, 
    6675, 
    6676, 
    6677, 
    6678, 
    6679, 
    6680, 
    6681, 
    6682, 
    6683, 
    6684, 
    6685, 
    6686, 
    6687, 
    6688, 
    6689, 
    6690, 
    6691, 
    6692, 
    6693, 
    6694, 
    6695, 
    6696, 
    6697, 
    6698, 
    6699, 
    6700, 
    6701, 
    6702, 
    6703, 
    6704, 
    6705, 
    6706, 
    6707, 
    6708 ;

 grid.vertices.xy =
  
    599996.822557256, 
    -1467643.50134789,
  
    617041.978149012, 
    -1488618.39186497,
  
    605475.42694971, 
    -1498596.3581024,
  
    637049.596036874, 
    -1535597.55748804,
  
    633428.937194709, 
    -1553981.79533051,
  
    617859.08859944, 
    -1564838.46280178,
  
    635152.111400938, 
    -1564944.12513423,
  
    642927.583637073, 
    -1580615.75725189,
  
    663884.775192954, 
    -1591957.22048923,
  
    653676.65921791, 
    -1603963.34948757,
  
    639909.27637197, 
    -1595860.34084325,
  
    623916.545439017, 
    -1581772.8788532,
  
    609287.440690019, 
    -1586024.9830141,
  
    617960.376662641, 
    -1603913.84687456,
  
    592366.922504426, 
    -1585293.32044808,
  
    575846.308110438, 
    -1595636.09454666,
  
    560656.978463049, 
    -1593603.70522026,
  
    557621.544813263, 
    -1608511.86053834,
  
    579062.083615133, 
    -1607670.02035482,
  
    597935.054741093, 
    -1619633.28461764,
  
    608426.603053189, 
    -1632557.08402587,
  
    622049.269193125, 
    -1639342.00023791,
  
    585626.269664076, 
    -1632812.53323796,
  
    567707.806383999, 
    -1637937.35139501,
  
    574285.875327318, 
    -1652373.02345297,
  
    539990.954595025, 
    -1660299.5805645,
  
    552158.341771438, 
    -1671266.4477982,
  
    561303.142055462, 
    -1659140.08332955,
  
    563469.662913299, 
    -1676920.77156953,
  
    549491.277327977, 
    -1682711.97478997,
  
    522644.166007665, 
    -1682385.13935785,
  
    538773.403941157, 
    -1691938.41283498,
  
    551453.508752352, 
    -1709878.50206845,
  
    538849.022836563, 
    -1699531.19681355,
  
    531332.293798802, 
    -1713784.27016222,
  
    515990.997857658, 
    -1723690.46546872,
  
    523794.121268221, 
    -1738890.48997814,
  
    530352.186554638, 
    -1723247.63179461,
  
    526956.631667406, 
    -1762876.74412017,
  
    547577.642906156, 
    -1755908.64189482,
  
    535992.115400584, 
    -1769536.11196382,
  
    544412.068290073, 
    -1783516.94710103,
  
    544888.992334661, 
    -1804654.69830603,
  
    557539.0949247, 
    -1786262.21931792,
  
    559087.140613298, 
    -1802094.30615534,
  
    571087.91684416, 
    -1813746.08159983,
  
    592443.135264714, 
    -1814545.76214463,
  
    573171.843075505, 
    -1821686.52368878,
  
    598752.109116622, 
    -1828813.25570523,
  
    607783.188755292, 
    -1845481.55883819,
  
    584196.575526136, 
    -1844895.96485629,
  
    593973.237609081, 
    -1856680.04804867,
  
    576659.121627548, 
    -1857174.74710965,
  
    591749.983317349, 
    -1867150.50702882,
  
    608466.08049765, 
    -1861680.25712302,
  
    595240.171046477, 
    -1870742.99432006,
  
    577708.984860965, 
    -1875216.03056097,
  
    558368.554993092, 
    -1876373.08990264,
  
    546243.612839137, 
    -1865170.41444854,
  
    530070.725316502, 
    -1868716.10813343,
  
    541971.949563896, 
    -1896869.98245738,
  
    530116.237023802, 
    -1906700.37318348,
  
    545832.886381693, 
    -1911893.18913634,
  
    553514.03999388, 
    -1894458.13200588,
  
    552531.63225754, 
    -1917467.87497491,
  
    568704.813312807, 
    -1923553.87190448,
  
    562724.110890284, 
    -1941806.99842189,
  
    547806.337857531, 
    -1943181.29296229,
  
    544035.249453809, 
    -1958884.48210933,
  
    581878.164244435, 
    -1967425.83896455,
  
    599038.945337894, 
    -1966659.37410222,
  
    588321.668854021, 
    -1980865.9880826,
  
    594969.962857498, 
    -1994364.04775437,
  
    608088.258128144, 
    -2005235.25318227,
  
    605869.441875131, 
    -2022672.09180794,
  
    589070.518176922, 
    -2031936.2102103,
  
    609505.218356586, 
    -2031943.70086778,
  
    596524.087784728, 
    -2046180.21701889,
  
    582830.371932584, 
    -2053178.2729508,
  
    565906.2182134, 
    -2053754.1798751,
  
    579569.286816216, 
    -2064981.456475,
  
    564082.217668593, 
    -2071556.7149834,
  
    583097.476053925, 
    -2065293.538901,
  
    577720.863317935, 
    -2082910.18261981,
  
    606072.743974427, 
    -2089119.41181569,
  
    606868.221525771, 
    -2105982.64745411,
  
    629401.2304931, 
    -2099596.41416048,
  
    642779.758726903, 
    -2091988.71370558,
  
    660263.411157939, 
    -2090224.82030986,
  
    673969.095951637, 
    -2097839.54355319,
  
    671043.639428084, 
    -2080257.05555026,
  
    680350.872047105, 
    -2064837.12915545,
  
    691822.31114363, 
    -2052866.61511691,
  
    703139.982951545, 
    -2063542.51564593,
  
    713667.839045186, 
    -2050306.71881543,
  
    718258.325161152, 
    -2033884.03154847,
  
    730862.091729434, 
    -2042411.19921909,
  
    740870.180187244, 
    -2029428.72616296,
  
    756654.103209579, 
    -2026564.84982025,
  
    820134.719334167, 
    -2019636.03860225,
  
    820720.862289284, 
    -2035562.01444615,
  
    801050.540466718, 
    -2043428.61254058,
  
    793464.073238673, 
    -2057061.42814829,
  
    807682.31871975, 
    -2047086.59871957,
  
    785337.519900088, 
    -2074206.75274134,
  
    801261.09179736, 
    -2083246.37560635,
  
    784943.404871501, 
    -2084687.30376716,
  
    768580.614002316, 
    -2100165.0560147,
  
    769620.276051351, 
    -2120234.26244811,
  
    764883.733473146, 
    -2135304.976327,
  
    761859.992231457, 
    -2120026.49267042,
  
    740883.582838011, 
    -2151196.95564317,
  
    756223.52968957, 
    -2141437.6531001,
  
    746512.951302371, 
    -2175515.3317263,
  
    749898.153309659, 
    -2191249.64009397,
  
    733030.922392994, 
    -2185280.78909307,
  
    716388.688497856, 
    -2185014.61091724,
  
    718860.960873025, 
    -2204197.71658402,
  
    704887.378833012, 
    -2216795.22819517,
  
    686225.452117889, 
    -2213862.1708261,
  
    685966.121587771, 
    -2232520.55232587,
  
    672412.841352911, 
    -2224815.18927339,
  
    660044.472208028, 
    -2271009.6079149,
  
    642791.455634702, 
    -2271078.03300933,
  
    628988.080822043, 
    -2264737.89756954,
  
    612413.085006836, 
    -2251370.71437407,
  
    602939.750367195, 
    -2269191.91576091,
  
    613229.324581892, 
    -2281847.71631581,
  
    597176.028608925, 
    -2286606.06493762,
  
    583864.50144181, 
    -2274548.31246043,
  
    580995.602712801, 
    -2298096.11713397,
  
    565317.21433193, 
    -2309866.99248609,
  
    546892.952606522, 
    -2316955.95154238,
  
    538510.827670892, 
    -2302894.91059202,
  
    524397.060310453, 
    -2296791.75979757,
  
    518618.999021773, 
    -2281311.97953864,
  
    499279.538017732, 
    -2272566.20012115,
  
    495399.510817439, 
    -2287915.60701035,
  
    479354.366601444, 
    -2291598.96936532,
  
    493902.842564206, 
    -2297354.90651581,
  
    496103.712388156, 
    -2313757.54451568,
  
    508897.972266014, 
    -2321991.95370718,
  
    517831.932361188, 
    -2336368.41102793,
  
    536399.362594251, 
    -2336957.79966529,
  
    537128.29078788, 
    -2352284.04451608,
  
    529701.615414277, 
    -2365600.79516326,
  
    517458.153278147, 
    -2374648.0966305,
  
    512990.982882853, 
    -2389123.29764135,
  
    496587.725527473, 
    -2390707.44675077,
  
    497287.241750833, 
    -2423320.06614865,
  
    482456.071124661, 
    -2433573.66203027,
  
    490076.545899562, 
    -2464898.43371563,
  
    478621.365026122, 
    -2475339.18664347,
  
    475650.996609472, 
    -2511498.78012441,
  
    460046.826137588, 
    -2511347.84949026,
  
    460736.191649256, 
    -2526832.63103416,
  
    464778.401857897, 
    -2542617.59731934,
  
    448735.460895958, 
    -2546616.33896791,
  
    438142.05227967, 
    -2560035.09182799,
  
    423944.517449276, 
    -2550713.77516639,
  
    407256.946645886, 
    -2557304.80103318,
  
    376506.503686136, 
    -2555558.37726139,
  
    345497.118341226, 
    -2564065.66118637,
  
    335537.523859917, 
    -2575942.16808307,
  
    327907.573777712, 
    -2558372.56275414,
  
    312918.891556072, 
    -2560031.94921798,
  
    302665.448533652, 
    -2571381.01483894,
  
    304489.841051073, 
    -2587086.99931238,
  
    316457.010824574, 
    -2596072.22837505,
  
    308628.186530785, 
    -2613997.52716879,
  
    299162.539835562, 
    -2625580.85415338,
  
    306256.423957815, 
    -2642250.25989801,
  
    292534.220322869, 
    -2651687.63997494,
  
    285112.236085715, 
    -2665810.85991478,
  
    273685.601612154, 
    -2651056.13107707,
  
    256169.760086419, 
    -2660931.82892899,
  
    246479.215008004, 
    -2673208.50119477,
  
    233932.894716745, 
    -2681850.53708253,
  
    240133.411083089, 
    -2696886.15235816,
  
    242115.827141507, 
    -2713846.37582108,
  
    233859.919207165, 
    -2730508.84699829,
  
    217018.776276819, 
    -2726153.90573435,
  
    185562.566131634, 
    -2724310.00212761,
  
    189444.799875338, 
    -2757600.0054743,
  
    199648.036208106, 
    -2771820.59612334,
  
    211948.853733267, 
    -2782512.893026,
  
    214420.222189228, 
    -2798924.09388864,
  
    222642.390642089, 
    -2814377.65334256,
  
    208152.160074673, 
    -2810276.03963643,
  
    196548.329594761, 
    -2822109.71338342,
  
    181825.079922124, 
    -2819303.81799116,
  
    169949.532115448, 
    -2830169.76358297,
  
    182366.604104938, 
    -2840578.89944124,
  
    197885.454078055, 
    -2848760.26280454,
  
    212612.485896848, 
    -2841768.22747355,
  
    220307.70677636, 
    -2872318.91152836,
  
    219066.016630954, 
    -2888977.30927261,
  
    203945.233760596, 
    -2891191.85475112,
  
    173870.582042455, 
    -2871475.87827476,
  
    161338.724179949, 
    -2882802.63143052,
  
    171530.595220742, 
    -2896140.2311469,
  
    144471.359365084, 
    -2914754.64808141,
  
    156111.344611211, 
    -2925405.46889947,
  
    161749.378270937, 
    -2940100.81562259,
  
    130160.258967119, 
    -2937160.17475881,
  
    133104.612740586, 
    -2953919.78250438,
  
    131274.750147069, 
    -2970277.58644077,
  
    119330.777533487, 
    -2981313.51602797,
  
    102921.652579148, 
    -2988174.49542961,
  
    97012.6190188243, 
    -3002963.66114355,
  
    96237.0101772401, 
    -3018579.6209029,
  
    114390.227676636, 
    -3017022.23727767,
  
    98816.2010290153, 
    -3022496.87748325,
  
    100643.98809369, 
    -3037656.8716466,
  
    118320.786289989, 
    -3042049.45885216,
  
    128708.565507661, 
    -3054324.65413796,
  
    143270.000198339, 
    -3064005.58362022,
  
    132441.510398911, 
    -3096052.67961959,
  
    148385.96010693, 
    -3088848.64965231,
  
    138985.941945303, 
    -3100555.33987659,
  
    143994.174196631, 
    -3116685.14582287,
  
    129168.555054379, 
    -3119536.8885624,
  
    116784.865314011, 
    -3111107.9809804,
  
    135961.089360004, 
    -3137655.94453302,
  
    115484.243260551, 
    -3134638.37850104,
  
    136734.714339118, 
    -3158315.8395043,
  
    125980.98608503, 
    -3168756.68045057,
  
    110770.259781252, 
    -3165865.85345473,
  
    95529.894619105, 
    -3170113.34953979,
  
    101346.479715687, 
    -3185001.88265003,
  
    84769.528677649, 
    -3184939.68441016,
  
    68817.8036693526, 
    -3188750.430923,
  
    77671.5954732234, 
    -3210245.06680907,
  
    79347.7593644123, 
    -3226339.7637256,
  
    62040.4726854371, 
    -3236121.72640818,
  
    57843.2932334531, 
    -3251028.73704847,
  
    45087.3737285164, 
    -3242080.00507345,
  
    40696.0400381137, 
    -3257835.33651406,
  
    26227.1953626771, 
    -3252299.52892412,
  
    31337.0701969618, 
    -3237129.06218311,
  
    14967.2287788721, 
    -3222589.97020655,
  
    6.74773582751912, 
    -3215439.96372668,
  
    -394.724310718557, 
    -3198496.87871648,
  
    14917.2065083381, 
    -3192058.13116043,
  
    10046.4872240646, 
    -3177107.10151919,
  
    -5262.83063883138, 
    -3178951.51580257,
  
    11008.9240686823, 
    -3155215.27102774,
  
    -5387.67624496139, 
    -3147224.85889749,
  
    -38599.5712505017, 
    -3166379.78296383,
  
    -53242.8702639006, 
    -3160913.71536094,
  
    -60847.793957181, 
    -3174087.10602726,
  
    -65269.5923670001, 
    -3191542.98754293,
  
    -80521.4509424735, 
    -3199335.76821522,
  
    -96937.557468546, 
    -3202758.02931014,
  
    -113615.320700585, 
    -3201929.71110913,
  
    -129573.617653779, 
    -3196193.79688479,
  
    -150139.454469544, 
    -3201956.80999578,
  
    -154647.669547014, 
    -3187532.9123752,
  
    -149553.122970107, 
    -3172324.39389477,
  
    -165552.438407602, 
    -3144787.0538492,
  
    -153800.851174817, 
    -3131734.38114436,
  
    -174116.353934781, 
    -3135860.50263413,
  
    -166468.551151571, 
    -3119568.50181418,
  
    -167546.931660124, 
    -3103939.84684524,
  
    -176733.015303117, 
    -3092109.00402053,
  
    -194808.472937464, 
    -3093371.6730061,
  
    -185493.621820441, 
    -3081248.47514137,
  
    -202524.689630037, 
    -3079001.8936546,
  
    -206554.270396721, 
    -3062655.72595214,
  
    -218878.701259655, 
    -3047329.73841277,
  
    -232822.499573229, 
    -3012848.99276036,
  
    -249980.143612989, 
    -3015681.63609802,
  
    -269139.236270634, 
    -3024793.71247331,
  
    -265520.244434425, 
    -3009997.86958332,
  
    -239278.936114116, 
    -2992297.35923381,
  
    -232971.677485853, 
    -2975753.64258289,
  
    -241566.784384337, 
    -2962320.37117608,
  
    -219324.765584111, 
    -2948890.57864396,
  
    -233070.072068933, 
    -2940968.81857824,
  
    -217464.436249718, 
    -2934512.63550296,
  
    -223014.503056476, 
    -2919120.47477954,
  
    -239114.138990726, 
    -2915591.0914407,
  
    -248876.681507542, 
    -2903840.09548442,
  
    -287501.060903448, 
    -2904069.32084971,
  
    -269050.840177648, 
    -2900501.0952945,
  
    -267831.653346559, 
    -2885070.31678875,
  
    -250306.436728422, 
    -2881720.5369205,
  
    -222806.028538612, 
    -2858118.1962359,
  
    -230121.042794647, 
    -2842733.05344117,
  
    -227051.463932704, 
    -2824909.70058985,
  
    -209703.960101086, 
    -2818448.54708609,
  
    -227190.345606308, 
    -2816133.81015574,
  
    -214354.739354206, 
    -2805052.69917265,
  
    -216868.664820979, 
    -2786261.64450335,
  
    -232922.869096315, 
    -2779780.16809149,
  
    -219679.202580755, 
    -2767348.05537136,
  
    -229560.873700721, 
    -2752250.83561551,
  
    -236155.938464656, 
    -2736001.91529863,
  
    -225874.595243235, 
    -2717865.0893613,
  
    -244901.150299487, 
    -2706900.05298834,
  
    -261610.04478603, 
    -2711321.95657997,
  
    -245966.690916981, 
    -2693847.27230657,
  
    -235965.912292405, 
    -2676850.17291292,
  
    -234653.799205924, 
    -2660698.29906732,
  
    -252298.381444636, 
    -2660910.38136035,
  
    -263052.529156504, 
    -2648779.29296776,
  
    -240323.724843729, 
    -2641370.46829219,
  
    -226882.17435601, 
    -2610640.13030017,
  
    -205391.740719998, 
    -2587693.02997633,
  
    -204100.624637902, 
    -2553726.26485768,
  
    -206413.395874118, 
    -2535217.66487078,
  
    -217325.842798356, 
    -2522593.03300008,
  
    -227020.987302788, 
    -2492036.41887495,
  
    -211100.414744561, 
    -2482073.62495913,
  
    -205278.429883298, 
    -2464775.67800222,
  
    -206379.010625999, 
    -2419638.25568673,
  
    -222254.693093645, 
    -2392782.61238131,
  
    -219457.883502379, 
    -2374714.93902128,
  
    -232816.115480039, 
    -2365017.66198651,
  
    -248455.544475579, 
    -2367878.86326918,
  
    -219284.683934888, 
    -2324943.81583152,
  
    -218211.430335375, 
    -2304292.37043055,
  
    -200578.125323671, 
    -2301155.0121495,
  
    -189049.462953933, 
    -2280050.67549737,
  
    -195276.9390892, 
    -2262769.50141518,
  
    -205074.183187056, 
    -2250008.0004881,
  
    -199054.518048628, 
    -2234731.22690111,
  
    -199093.886172423, 
    -2202283.24362502,
  
    -206219.338454788, 
    -2188447.72098008,
  
    -194726.992507607, 
    -2175880.86346619,
  
    -203014.888538795, 
    -2135945.28757559,
  
    -200893.929973518, 
    -2118219.82645559,
  
    -207245.670140676, 
    -2103462.19600971,
  
    -202967.245200415, 
    -2088865.52861799,
  
    -211003.601486829, 
    -2071566.25792451,
  
    -211071.433925953, 
    -2055998.99185541,
  
    -221657.612807446, 
    -2043785.17632004,
  
    -220340.908227363, 
    -2028243.9332106,
  
    -226291.855956512, 
    -2011953.4937414,
  
    -225315.00496974, 
    -1997005.03562934,
  
    -217749.132319199, 
    -1983940.5288894,
  
    -249415.971701471, 
    -1977808.58698441,
  
    -238316.793848619, 
    -1964518.0007311,
  
    -254594.427300835, 
    -1980232.04100681,
  
    -255760.038406089, 
    -1946887.50151748,
  
    -246625.937197696, 
    -1934133.1021162,
  
    -261064.58460049, 
    -1948491.42751938,
  
    -252021.63246975, 
    -1927457.73264072,
  
    -267216.931055371, 
    -1938270.70243404,
  
    -278540.24052946, 
    -1905275.74368816,
  
    -265479.85112598, 
    -1897348.55902353,
  
    -280562.651430265, 
    -1896926.63214665,
  
    -303606.803696643, 
    -1848455.92838106,
  
    -303782.529114953, 
    -1832783.99103054,
  
    -322320.536635711, 
    -1806901.04927511,
  
    -317466.666844074, 
    -1791756.73024655,
  
    -328174.551531031, 
    -1762344.16604961,
  
    -319557.793145059, 
    -1749731.20192065,
  
    -326862.296007619, 
    -1735167.33498215,
  
    -326257.342548323, 
    -1720007.32330928,
  
    -330487.451009677, 
    -1703845.92547916,
  
    -331660.72938743, 
    -1688296.99375894,
  
    -329559.107929866, 
    -1673271.99397757,
  
    -322606.63999224, 
    -1656012.82896668,
  
    -331603.262595395, 
    -1643996.77441698,
  
    -333244.706898518, 
    -1625651.90612371,
  
    -347449.104443163, 
    -1598856.0529311,
  
    -361966.985712115, 
    -1590839.47377938,
  
    -360656.712227769, 
    -1574312.60771227,
  
    -364799.913790544, 
    -1558760.56009748,
  
    -356054.542411412, 
    -1545754.70067938,
  
    -343722.064654382, 
    -1534317.7456381,
  
    -359979.453749701, 
    -1531162.1409039,
  
    -358271.175186661, 
    -1514819.16752519,
  
    -373741.571388615, 
    -1509522.83777256,
  
    -375578.695947983, 
    -1493828.60361557,
  
    -382547.051292464, 
    -1479254.58994222,
  
    -392419.765990139, 
    -1467929.74789729,
  
    -407852.620826452, 
    -1465182.92081781,
  
    -405216.056937495, 
    -1448380.66123113,
  
    -415496.727098011, 
    -1436104.93294652,
  
    -432511.185369504, 
    -1437111.08617349,
  
    -435705.436652655, 
    -1422300.42907999,
  
    -453048.8328734, 
    -1421807.48106649,
  
    -456974.476482074, 
    -1404657.32026767,
  
    -472402.728442764, 
    -1405808.80712945,
  
    -478853.203569341, 
    -1421389.39874681,
  
    -487029.91800206, 
    -1408653.34632007,
  
    -501998.023392359, 
    -1406837.15346365,
  
    -529051.877679414, 
    -1425362.84153104,
  
    -533728.235721044, 
    -1411147.79886936,
  
    -520457.122103705, 
    -1403691.11927057,
  
    -529161.392157512, 
    -1389621.06773091,
  
    -542400.742001857, 
    -1397836.17852411,
  
    -551217.614302659, 
    -1409947.23789071,
  
    -551092.124459481, 
    -1393301.49485877,
  
    -564842.689982711, 
    -1384083.20819803,
  
    -566192.690705608, 
    -1400003.38720573,
  
    -589775.301238753, 
    -1397223.29736954,
  
    -594018.650428097, 
    -1380870.25801184,
  
    -606643.758217776, 
    -1369720.33388244,
  
    -591995.62554031, 
    -1365445.65145009,
  
    -580593.380954737, 
    -1351731.85516052,
  
    -563534.556613671, 
    -1356473.432509,
  
    -548097.826909387, 
    -1356312.71989514,
  
    -546245.53385827, 
    -1340582.5666354,
  
    -519823.692308829, 
    -1322774.9524882,
  
    -509263.856498909, 
    -1311091.50516966,
  
    -493138.770065682, 
    -1315644.14739789,
  
    -502153.173686184, 
    -1300953.84802769,
  
    -480681.977860791, 
    -1288113.35560483,
  
    -488532.603900899, 
    -1272525.96309518,
  
    -465001.745206455, 
    -1269816.53267053,
  
    -485868.522889535, 
    -1255070.08146643,
  
    -491071.469685074, 
    -1240675.48559922,
  
    -508577.63652049, 
    -1238693.02726031,
  
    -520666.90321914, 
    -1247992.1818737,
  
    -530413.481089036, 
    -1233518.98872825,
  
    -544062.277477091, 
    -1223445.08039853,
  
    -546894.889075033, 
    -1208104.72838778,
  
    -557514.686231328, 
    -1197437.81136034,
  
    -566705.873245934, 
    -1183561.61236553,
  
    -581999.095860129, 
    -1180826.20290492,
  
    -593994.283953859, 
    -1168912.57024886,
  
    -597210.185088166, 
    -1151006.05060057,
  
    -585473.733054595, 
    -1138741.38522315,
  
    -568624.119468542, 
    -1134164.46109178,
  
    -549049.939270905, 
    -1142460.3766678,
  
    -538028.497578035, 
    -1155646.77423591,
  
    -520761.17879946, 
    -1163260.29299992,
  
    -501252.578921299, 
    -1153211.98885815,
  
    -460321.971359158, 
    -1150858.56553846,
  
    -457992.394074483, 
    -1133369.89923009,
  
    -439295.514379038, 
    -1125314.99310818,
  
    -426307.975023091, 
    -1115000.89845595,
  
    -420154.588556536, 
    -1101321.29613533,
  
    -374323.263877425, 
    -1063332.15694111,
  
    -367380.284414047, 
    -1048251.89042273,
  
    -357045.95910033, 
    -1036822.5550876,
  
    -322668.685599335, 
    -1043236.68167264,
  
    -320867.280011626, 
    -1028375.11188286,
  
    -315952.611203316, 
    -1045211.98344634,
  
    -298956.599033367, 
    -1051611.52618077,
  
    -283621.667597959, 
    -1039879.02501008,
  
    -268429.933985319, 
    -1033360.11395522,
  
    -268024.601554565, 
    -1017457.25726107,
  
    -280793.988261146, 
    -1025837.54061011,
  
    -269862.73106157, 
    -1015389.28864996,
  
    -281981.241039186, 
    -988942.490572329,
  
    -286279.418900018, 
    -969395.059888699,
  
    -287170.902781069, 
    -929252.033513142,
  
    -276244.1295215, 
    -917684.385277408,
  
    -260386.639347146, 
    -916404.513668977,
  
    -246520.368644412, 
    -904631.453605587,
  
    -232656.097568701, 
    -916021.57733379,
  
    -215990.863609273, 
    -916417.817404604,
  
    -195081.480316733, 
    -939730.115786867,
  
    -179571.636382229, 
    -943520.346093975,
  
    -164869.934945163, 
    -939737.54253362,
  
    -148464.762651869, 
    -922077.991163736,
  
    -158337.619662624, 
    -910804.868627071,
  
    -143384.342852576, 
    -916807.344111395,
  
    -148571.516320375, 
    -932114.953404639,
  
    -142534.540022014, 
    -946896.4035838,
  
    -123179.895397576, 
    -947513.832536762,
  
    -105809.773549842, 
    -954291.812372389,
  
    -91535.7515399948, 
    -949626.669332604,
  
    -89662.2091306806, 
    -932564.012165232,
  
    -92502.7932239315, 
    -900250.565455638,
  
    -88405.0477086913, 
    -885185.732598869,
  
    -77700.0098145027, 
    -904424.878331874,
  
    -78251.1663895482, 
    -923197.042503439,
  
    -70720.2630032935, 
    -945641.080819456,
  
    -52503.9511522614, 
    -943510.138955465,
  
    -41018.8682136193, 
    -929627.82206615,
  
    -16092.589101121, 
    -931223.733754896,
  
    -16251.9336120708, 
    -913382.745854754,
  
    -3619.16739467235, 
    -901799.157816293,
  
    13810.0657845348, 
    -899417.298608448,
  
    -1101.07757978245, 
    -896982.60359058,
  
    -11153.3524399593, 
    -885892.066482085,
  
    4297.08762526923, 
    -891373.499805196,
  
    27418.4241023628, 
    -864603.181730471,
  
    47105.9194624623, 
    -869444.993631578,
  
    35793.6472625055, 
    -859200.441741757,
  
    48534.8014502257, 
    -848238.025993782,
  
    63662.8805470947, 
    -849020.24758928,
  
    49845.8934400715, 
    -833979.077390462,
  
    68492.1020225156, 
    -834167.821575196,
  
    74061.0763637313, 
    -848107.506555565,
  
    87095.0470467948, 
    -862518.21771608,
  
    91769.7241762524, 
    -847119.067115116,
  
    101735.846826675, 
    -858605.407808468,
  
    118967.094475927, 
    -861537.22930259,
  
    127265.839846432, 
    -876659.470068786,
  
    146102.91440922, 
    -862841.462746442,
  
    136922.425920445, 
    -877138.674388706,
  
    151591.050247843, 
    -881772.841918356,
  
    168435.866073579, 
    -872043.865559617,
  
    184764.742410385, 
    -870337.636279335,
  
    169011.545968815, 
    -877366.664382385,
  
    162145.193616233, 
    -890688.101919159,
  
    166816.464981168, 
    -910468.03752964,
  
    180770.894844903, 
    -904385.912975984,
  
    201403.34653577, 
    -881807.290454283,
  
    226880.663087271, 
    -910375.11921288,
  
    245765.754781322, 
    -907029.992997017,
  
    259689.933597989, 
    -898121.459262997,
  
    274806.006217963, 
    -882907.254000453,
  
    269977.469675481, 
    -903901.320538632,
  
    259652.549651027, 
    -916756.159643229,
  
    274473.775417502, 
    -925053.751527212,
  
    293308.644780176, 
    -928802.298647275,
  
    278428.471128816, 
    -940478.830837066,
  
    290029.378774525, 
    -951241.131096904,
  
    303651.757948012, 
    -958694.310664704,
  
    314742.552266049, 
    -973835.073208784,
  
    332164.401246034, 
    -974887.23698531,
  
    344168.170393331, 
    -986643.169859189,
  
    338411.853043953, 
    -1001756.07717071,
  
    353580.73458045, 
    -999038.476328637,
  
    368722.110569719, 
    -1002333.78169743,
  
    382164.123995248, 
    -1017287.23108434,
  
    391782.967900245, 
    -1035221.8086139,
  
    408673.947024964, 
    -1049898.52848852,
  
    422990.621204186, 
    -1056662.16060043,
  
    435712.674928821, 
    -1047805.89285091,
  
    455465.192215173, 
    -1022455.83784062,
  
    461272.430678037, 
    -1006243.9865846,
  
    477963.629796283, 
    -1009110.08124661,
  
    488298.601668349, 
    -1021453.36960119,
  
    487480.652661398, 
    -1036424.06862334,
  
    462337.676538163, 
    -1057603.56239036,
  
    453722.098816237, 
    -1072657.25259443,
  
    469274.378904715, 
    -1080426.63605024,
  
    484837.153115558, 
    -1083239.72934144,
  
    501560.296976321, 
    -1077475.61878795,
  
    512611.484771493, 
    -1066807.52984255,
  
    522333.8509203, 
    -1082446.99471411,
  
    522785.605415423, 
    -1102141.06510695,
  
    509071.120199388, 
    -1094557.11641383,
  
    489486.756303238, 
    -1118674.87004789,
  
    483138.242960074, 
    -1132336.00900571,
  
    478968.186056405, 
    -1149661.46899079,
  
    495064.19100172, 
    -1137629.90141019,
  
    508242.631750554, 
    -1169542.31225224,
  
    506683.599148506, 
    -1188269.52032417,
  
    508741.835653422, 
    -1209847.72705556,
  
    520933.715000832, 
    -1222584.23855928,
  
    516720.506253864, 
    -1239310.43668471,
  
    529487.006258496, 
    -1247442.86245844,
  
    539233.606757063, 
    -1260309.09308051,
  
    543334.797973156, 
    -1277859.22415745,
  
    551422.203635026, 
    -1293830.71225971,
  
    558716.194034449, 
    -1330049.82815952,
  
    557428.445980087, 
    -1345734.95846521,
  
    515100.684062406, 
    -1299770.11687941,
  
    498761.06153174, 
    -1289613.36134753,
  
    509794.509561259, 
    -1303853.2536537,
  
    492788.340387179, 
    -1294287.46566187,
  
    492435.134885253, 
    -1310390.32115756,
  
    479708.501391114, 
    -1331475.19598371,
  
    508150.649386576, 
    -1313048.28505897,
  
    484057.803200466, 
    -1342016.29231709,
  
    498149.148973091, 
    -1334109.16301402,
  
    509516.325107399, 
    -1354806.01220386,
  
    528077.835265022, 
    -1346723.75529379,
  
    515893.877948653, 
    -1360359.76875984,
  
    501983.01005663, 
    -1354160.11584207,
  
    486829.816718809, 
    -1351203.6201057,
  
    476920.691268503, 
    -1366132.02224636,
  
    493114.152968294, 
    -1365329.15242582,
  
    499414.141251299, 
    -1379126.70522071,
  
    486223.881839599, 
    -1394963.25929916,
  
    500909.446727018, 
    -1399722.42477841,
  
    515581.432806891, 
    -1391279.01378042,
  
    529508.244057617, 
    -1378801.48986119,
  
    542769.268960761, 
    -1351199.44416603,
  
    561905.407611796, 
    -1350467.48685763,
  
    564887.312043059, 
    -1370913.98233815,
  
    578203.108962924, 
    -1381075.24652397,
  
    573717.779004081, 
    -1397424.90873184,
  
    587820.491325503, 
    -1389017.91437879,
  
    585282.449391145, 
    -1409115.4190831,
  
    579181.138592149, 
    -1427028.92073017,
  
    589850.579808121, 
    -1439534.06389141,
  
    616570.186886932, 
    -1509689.88126534,
  
    626652.846039032, 
    -1522023.72327435,
  
    606032.781256749, 
    -1593607.59950528,
  
    603334.940076054, 
    -1637529.18301242,
  
    556880.419072166, 
    -1656247.87913007,
  
    529315.643778826, 
    -1742794.11819758,
  
    536414.736519547, 
    -1882703.44677765,
  
    562966.94572466, 
    -1964044.4600456,
  
    772898.511166779, 
    -2027094.27308182,
  
    789162.449240106, 
    -2026249.95549544,
  
    804880.100303007, 
    -2023546.47860933,
  
    797199.578435137, 
    -2060637.0712641,
  
    752109.068853679, 
    -2134874.94645744,
  
    750317.4041714, 
    -2158448.46514711,
  
    668386.190753031, 
    -2239876.07455229,
  
    665331.429477525, 
    -2255395.40860316,
  
    496098.252527416, 
    -2406559.50821892,
  
    486572.954902473, 
    -2449638.73092195,
  
    476027.797846604, 
    -2492803.46358963,
  
    391828.157943275, 
    -2556266.58133864,
  
    360442.439038996, 
    -2558690.20113426,
  
    201098.265254358, 
    -2725475.7698007,
  
    188717.529374784, 
    -2740313.5196081,
  
    216589.708014552, 
    -2856774.52021845,
  
    188607.827331905, 
    -2881503.21377366,
  
    158429.44641646, 
    -2906045.51493858,
  
    146229.790254538, 
    -2938921.68496978,
  
    136803.953174755, 
    -3079870.88469285,
  
    126530.928228571, 
    -3123843.79193645,
  
    125626.916176077, 
    -3147730.9848004,
  
    -21817.0554301363, 
    -3156405.71855461,
  
    -158129.219541569, 
    -3158920.37315059,
  
    -226492.777297361, 
    -3029681.97886978,
  
    -253230.46157584, 
    -3000171.88646825,
  
    -267318.885259677, 
    -2905311.30522561,
  
    -237487.159019663, 
    -2869479.75592582,
  
    -233019.793723756, 
    -2625713.37537766,
  
    -215163.128555407, 
    -2599610.02528434,
  
    -205461.438557792, 
    -2571445.19674932,
  
    -220991.501864246, 
    -2507098.03209536,
  
    -205728.464824518, 
    -2442417.04026413,
  
    -214831.039847277, 
    -2405757.9663566,
  
    -238009.419861855, 
    -2355278.07942935,
  
    -229448.533935436, 
    -2340453.90415072,
  
    -198041.326673477, 
    -2218556.82417678,
  
    -200341.826975075, 
    -2157018.54217017,
  
    -233117.307651455, 
    -1979618.97798968,
  
    -255408.909309467, 
    -1963172.55803401,
  
    -272061.323749362, 
    -1920489.00456313,
  
    -289004.542079257, 
    -1881853.96057842,
  
    -297322.454862021, 
    -1865119.56806078,
  
    -312678.418556357, 
    -1819625.2439672,
  
    -323211.498153224, 
    -1776983.4172181,
  
    -340602.386439145, 
    -1612118.39365105,
  
    -514997.741992544, 
    -1417032.44302069,
  
    -532800.007231137, 
    -1331611.08105654,
  
    -479231.921301301, 
    -1150480.58597047,
  
    -406283.417290555, 
    -1090634.60874536,
  
    -390402.976861883, 
    -1078108.78601342,
  
    -340286.528094795, 
    -1039226.90293715,
  
    -285929.810295058, 
    -948518.81100952,
  
    -206291.912263743, 
    -928802.815041984,
  
    -91796.3858164405, 
    -916263.510673397,
  
    15006.4949870762, 
    -878133.788810929,
  
    191571.347105092, 
    -894258.176291619,
  
    213872.85064684, 
    -896144.25307884,
  
    445730.547731789, 
    -1035385.83286506,
  
    474179.748274093, 
    -1045778.50197234,
  
    499567.027221062, 
    -1106850.05335804,
  
    500649.896021221, 
    -1154280.48444153,
  
    556329.874767618, 
    -1312777.32884163,
  
    544219.237338874, 
    -1330770.76748069,
  
    530071.52627525, 
    -1314741.94441543,
  
    494501.916025522, 
    -1321420.96561642,
  
    497313.39402048, 
    -1328034.25640048,
  
    536118.184248433, 
    -1365043.28696799,
  
    595261.888977816, 
    -1453194.88391859,
  
    -304163.439089111, 
    -1733927.30013996,
  
    1795.93283863856, 
    -2053236.0202706,
  
    169234.749774023, 
    -2724054.2382063,
  
    24682.5499358368, 
    -889630.091502159,
  
    750115.990062744, 
    -2108729.69788818,
  
    261498.356200842, 
    -930591.715025142,
  
    -8629.51983237093, 
    -2754204.59831192,
  
    -349287.05244756, 
    -1466673.26369644,
  
    13110.4491987698, 
    -2485066.6029544,
  
    -253682.433854771, 
    -1351650.19779157,
  
    -396402.75649863, 
    -1415472.10341761,
  
    55922.5982228134, 
    -3146369.31737758,
  
    434644.061163753, 
    -1916560.81913983,
  
    30022.5168724418, 
    -2883634.12440829,
  
    111217.816668445, 
    -1062857.82646478,
  
    -272643.590276208, 
    -931814.63321008,
  
    40310.5151585222, 
    -2216229.25037406,
  
    -341293.288076063, 
    -1518157.82359789,
  
    188740.60852598, 
    -2666801.75734237,
  
    516952.99414747, 
    -2217745.4326671,
  
    -196006.368503094, 
    -1504044.31747529,
  
    509817.18371937, 
    -2256250.3698005,
  
    -202511.75408984, 
    -2340649.4273344,
  
    195235.752033628, 
    -906264.758035299,
  
    348066.577963366, 
    -1418160.9642862,
  
    330244.252120556, 
    -1764967.02221468,
  
    392302.778790871, 
    -2506373.02175304,
  
    -213373.564641972, 
    -2638418.89350739,
  
    82515.6859318957, 
    -2920518.34094367,
  
    93842.4729286787, 
    -1935930.35455362,
  
    55154.6041994403, 
    -2165559.46658803,
  
    208760.858695465, 
    -2547560.29638038,
  
    -147154.230363912, 
    -2280774.51843205,
  
    -538986.166189915, 
    -1194533.66417591,
  
    -81981.5474117332, 
    -2339769.60370752,
  
    533382.658580032, 
    -1520816.42332708,
  
    6835.99196982471, 
    -3032329.70601798,
  
    -373294.689449011, 
    -1431920.1304902,
  
    -315931.332954023, 
    -1060060.73175432,
  
    -271054.179528008, 
    -1657621.29592591,
  
    -337689.086281315, 
    -1569087.77046953,
  
    544244.755058013, 
    -1385009.29769172,
  
    35471.9483733586, 
    -2976877.26320878,
  
    446655.094860524, 
    -1304791.76599469,
  
    225578.02204359, 
    -2014297.15381669,
  
    -61581.0761298485, 
    -2720438.64972053,
  
    -201786.211471, 
    -965980.289482921,
  
    -56536.808472772, 
    -2155013.03180094,
  
    533816.625679814, 
    -2011448.44795036,
  
    -181733.392384906, 
    -2790249.88472099,
  
    -310355.846717519, 
    -1258041.00764588,
  
    226634.885701058, 
    -2548716.81125921,
  
    -154306.538117493, 
    -1150041.73529562,
  
    -31969.4420077212, 
    -2823935.82757801,
  
    122746.713755373, 
    -3082716.31788367,
  
    -153738.169718258, 
    -2948383.69036657,
  
    65300.0983651161, 
    -3074179.53527113,
  
    -10036.1581591176, 
    -977410.750738761,
  
    -177938.600541415, 
    -2178762.89367945,
  
    412000.93107409, 
    -1715298.12099847,
  
    373508.901428734, 
    -1945615.99722148,
  
    526399.267035389, 
    -2169421.12463473,
  
    -481084.007476912, 
    -1345315.20624712,
  
    123560.96119428, 
    -1455857.23149751,
  
    118517.805400607, 
    -1812016.77671432,
  
    479734.381719668, 
    -2308993.48410755,
  
    529603.659245672, 
    -1852841.8798663,
  
    -127212.743487621, 
    -2847262.01520902,
  
    -108692.071898878, 
    -1967136.96845261,
  
    646613.789891668, 
    -2149706.96874034,
  
    -154569.398573585, 
    -2103245.6433832,
  
    -21816.7402028842, 
    -2489069.81636013,
  
    111877.631683554, 
    -2285249.9208371,
  
    -139957.421596598, 
    -3183788.32618935,
  
    117682.700590506, 
    -2624395.29234748,
  
    500802.332512337, 
    -1510013.59876383,
  
    712799.029612396, 
    -2128802.41841667,
  
    651435.942475206, 
    -2243356.97984559,
  
    -459181.947490471, 
    -1246531.24171248,
  
    394997.904825725, 
    -2427652.03351674,
  
    -176593.974020207, 
    -1608887.32884925,
  
    -125300.517003899, 
    -1900653.59395196,
  
    -50707.8918102365, 
    -2904768.27834328,
  
    231807.954783585, 
    -1131349.46567631,
  
    455574.906669408, 
    -1974276.89102604,
  
    -148481.681890453, 
    -2759786.63856107,
  
    151634.113364083, 
    -2208070.85743955,
  
    491640.349980239, 
    -2228400.62065778,
  
    40143.5489017021, 
    -2815435.35964929,
  
    -271424.643700431, 
    -1049408.74939827,
  
    175175.829930173, 
    -2495846.20252054,
  
    -476317.965570629, 
    -1309566.45826041,
  
    50448.1628971147, 
    -2992828.153552,
  
    173990.944471545, 
    -1124313.39610655,
  
    86074.5401532858, 
    -3031444.14621551,
  
    186689.1211911, 
    -1697114.70415638,
  
    169919.367563909, 
    -1996206.3041275,
  
    -33412.1430990551, 
    -2603652.43921135,
  
    304817.458358714, 
    -1798591.54438949,
  
    -94448.9825616807, 
    -1492462.82533237,
  
    -84661.3862814889, 
    -1857167.163756,
  
    376512.367024302, 
    -2472755.1948808,
  
    149453.335521868, 
    -909214.004566437,
  
    456261.692186236, 
    -1252474.2935959,
  
    675646.862229071, 
    -2113721.84223907,
  
    -232508.079546835, 
    -2886557.8349448,
  
    346096.397620723, 
    -2289296.61732116,
  
    -448841.33537553, 
    -1353929.60120132,
  
    -86725.0729121761, 
    -2523369.23688906,
  
    362030.703797544, 
    -1389678.02480503,
  
    -224078.982482562, 
    -1011796.03243022,
  
    629013.067051341, 
    -2244023.66548672,
  
    34313.2143763486, 
    -1540817.15997679,
  
    100018.124002993, 
    -1838477.36041525,
  
    -214206.643996819, 
    -2885789.74036668,
  
    16960.8147084143, 
    -957907.165359126,
  
    552155.977363301, 
    -2144721.14861874,
  
    73002.9783848179, 
    -2736264.2138397,
  
    -446269.626561783, 
    -1332738.11870293,
  
    354508.554431377, 
    -2259778.73741402,
  
    -186619.951858043, 
    -2468691.65122514,
  
    43830.646951843, 
    -3221002.8541427,
  
    -30534.1173792042, 
    -2373967.55708878,
  
    -182970.518446574, 
    -1142408.33292682,
  
    295351.928387137, 
    -2601051.95187579,
  
    -319585.884100033, 
    -1233243.84634487,
  
    389035.953704793, 
    -1678216.48786734,
  
    353481.333480503, 
    -1267594.53588915,
  
    -334296.005811032, 
    -1061851.38047133,
  
    -112504.776179752, 
    -3074807.97493699,
  
    -35269.4835285701, 
    -1679201.89969485,
  
    -40743.7020283927, 
    -2048554.32659815,
  
    255114.794082602, 
    -957442.387488828,
  
    173738.614400098, 
    -2664243.78397846,
  
    100157.006282778, 
    -1871182.49696506,
  
    187443.810987886, 
    -2773803.82137115,
  
    -310485.654404034, 
    -1528737.09134397,
  
    561440.048592836, 
    -2276872.94112061,
  
    704180.108003747, 
    -2112158.4264316,
  
    617409.466253902, 
    -1545600.35539174,
  
    510236.866847709, 
    -1429989.99226947,
  
    100491.4481213, 
    -1951072.3791222,
  
    -15621.2789383131, 
    -2983710.60537153,
  
    382708.113442698, 
    -2275007.91502095,
  
    -290288.939924713, 
    -1178799.42802415,
  
    -140726.394893563, 
    -2557091.07312841,
  
    479047.045173522, 
    -1169028.79714946,
  
    148663.587009856, 
    -1433406.31217889,
  
    -337435.650945065, 
    -1589118.24359689,
  
    -555263.683635115, 
    -1156925.34582068,
  
    -137473.161885122, 
    -2582893.92154249,
  
    251025.034860599, 
    -1470873.54940047,
  
    325336.762555004, 
    -1776301.12713584,
  
    69724.2512552104, 
    -2683830.90078616,
  
    44026.6863822615, 
    -943185.090678578,
  
    421013.662903728, 
    -1885519.67128756,
  
    -308742.204835917, 
    -1779254.67446722,
  
    385683.461069757, 
    -2263767.19043894,
  
    45889.387794272, 
    -2517489.8304139,
  
    -486682.284285689, 
    -1207238.20683588,
  
    78050.6103837294, 
    -3067288.59413224,
  
    245041.778099419, 
    -2522172.35352962,
  
    -266561.323310545, 
    -1346201.22932402,
  
    -28545.7112074226, 
    -3037756.91414264,
  
    -302538.944698617, 
    -1069938.55707754,
  
    -39348.6614890479, 
    -3138159.68766861,
  
    117525.512105695, 
    -1669745.20559944,
  
    487685.532183341, 
    -1240887.29538204,
  
    -524492.543119313, 
    -1356198.01248917,
  
    -21143.8769798656, 
    -3142156.63737706,
  
    -254997.898918288, 
    -1661469.08220864,
  
    -134712.852499614, 
    -2076989.02703052,
  
    459898.049990963, 
    -1091494.7999495,
  
    -98143.3350585993, 
    -1941517.58547446,
  
    121957.939433765, 
    -2734101.51834742,
  
    -105699.684252385, 
    -3153650.98754832,
  
    -130705.766442595, 
    -2442195.94660628,
  
    -313708.854332955, 
    -1473428.56392247,
  
    -360569.434920236, 
    -1281671.72088767,
  
    579864.883870043, 
    -1552886.27184766,
  
    307347.828497626, 
    -1929708.07940286,
  
    -105103.073766216, 
    -2846891.25204594,
  
    235069.103236786, 
    -1153141.26989539,
  
    -203783.443889156, 
    -3009693.04036093,
  
    173307.899571936, 
    -2239060.62733401,
  
    -321863.058923012, 
    -1388878.43467301,
  
    66556.9485237935, 
    -2626115.27769872,
  
    448391.035804795, 
    -1207334.66519172,
  
    -64703.5295198509, 
    -1477134.60200837,
  
    595878.642817801, 
    -2122998.21846382,
  
    -251752.19864697, 
    -951873.105838502,
  
    469423.962484988, 
    -1400385.42292464,
  
    465332.792928619, 
    -1734947.70860432,
  
    418769.556837988, 
    -2533192.27019981,
  
    -118513.007920875, 
    -2618052.35969358,
  
    275650.241956499, 
    -989269.002775698,
  
    218479.118076112, 
    -1916726.28518752,
  
    390000.937054164, 
    -1122140.44787373,
  
    182729.833939054, 
    -2203465.00153638,
  
    256635.35398127, 
    -2561720.39524835,
  
    552922.884708851, 
    -1997436.38275034,
  
    51096.2004251115, 
    -2413995.94954501,
  
    -347622.951281408, 
    -1300585.26135613,
  
    -395797.615027426, 
    -1178873.26605876,
  
    -129945.526180617, 
    -1662023.96868142,
  
    545382.061698732, 
    -1826681.92401964,
  
    -99427.4580976928, 
    -2954282.79569588,
  
    -286269.948828412, 
    -1809519.48524884,
  
    87113.9230291106, 
    -2038390.39080303,
  
    85544.2151224723, 
    -2722743.27585476,
  
    -217480.051760831, 
    -975207.59423318,
  
    -184854.252087385, 
    -2122307.96112562,
  
    198705.608786915, 
    -919042.550656651,
  
    -93836.6670847514, 
    -2767321.67728997,
  
    -334313.511006956, 
    -1386430.08840195,
  
    98161.9171697247, 
    -2510419.87648155,
  
    -216165.920700221, 
    -1275538.71644006,
  
    -173697.368292189, 
    -2819560.19669682,
  
    105164.403219364, 
    -3152985.05619297,
  
    514204.206676787, 
    -1908343.78239595,
  
    111955.2188436, 
    -2905912.97542482,
  
    36139.9674095206, 
    -1008128.59047921,
  
    -43631.452716633, 
    -2201819.11397912,
  
    503406.686756513, 
    -2373265.71132885,
  
    498794.767885969, 
    -1914483.49919246,
  
    546408.759637186, 
    -2126377.48550397,
  
    -278070.646307848, 
    -1520862.8893832,
  
    -124682.909313433, 
    -3125305.04975323,
  
    261718.263384154, 
    -1432659.52807132,
  
    248498.366294181, 
    -1783132.55544706,
  
    456697.988119055, 
    -2454373.47914467,
  
    3108.06933450172, 
    -2892781.94709363,
  
    15944.5732484779, 
    -1947932.89908692,
  
    509565.371982183, 
    -1274784.75007165,
  
    -25508.4750525022, 
    -2141592.61221496,
  
    124633.097674657, 
    -2526219.65882899,
  
    -44363.0477890104, 
    -2282550.48427915,
  
    268299.170211709, 
    -2626615.77671173,
  
    -170927.744564671, 
    -2290158.36841542,
  
    504506.703387049, 
    -1443754.83647001,
  
    81983.1791673189, 
    -3007858.00259505,
  
    446403.091170249, 
    -2520331.5961555,
  
    -396455.768916185, 
    -1100141.91140754,
  
    329334.693294069, 
    -2533555.96816614,
  
    -306383.01063807, 
    -1650776.66271526,
  
    517637.882063997, 
    -2356241.58715062,
  
    72195.7433644753, 
    -2971493.25269806,
  
    364021.579634997, 
    -1238083.18892928,
  
    314038.362264458, 
    -1998904.74486233,
  
    -162204.183862086, 
    -2718862.44904005,
  
    23661.5903783537, 
    -2175453.70102061,
  
    517148.489610721, 
    -2097188.31601691,
  
    -94624.6810698781, 
    -2800137.68282333,
  
    288832.191843747, 
    -2563185.11446934,
  
    -115151.696963708, 
    -1070606.50767475,
  
    53521.2547609419, 
    -2826575.22148907,
  
    482867.817690761, 
    -1106149.74000654,
  
    -74080.3351446473, 
    -2965722.51028961,
  
    6393.61955462222, 
    -3135050.63933461,
  
    60743.4964701253, 
    -1033911.76782989,
  
    -498342.95643551, 
    -1178207.88701371,
  
    325342.543770807, 
    -1708304.49882823,
  
    295205.234021157, 
    -1965073.80609896,
  
    496599.791796643, 
    -2246811.77992632,
  
    -169437.067603331, 
    -2563865.31519191,
  
    434466.650713208, 
    -1752606.31354479,
  
    38496.6603070867, 
    -1470140.20004472,
  
    40146.9240442806, 
    -1829432.31829879,
  
    440129.016917491, 
    -2360694.44042912,
  
    -186589.971578988, 
    -1979139.51298559,
  
    633387.258110873, 
    -2154061.72410129,
  
    743661.200623092, 
    -2049881.62956031,
  
    -121543.34552556, 
    -2463772.23089953,
  
    204817.222892284, 
    -2286855.67785758,
  
    -461169.212904675, 
    -1334194.8195835,
  
    41327.7487904334, 
    -2586657.7876226,
  
    514110.458867637, 
    -1615038.77663987,
  
    -185415.398267792, 
    -976346.552208117,
  
    528186.330238475, 
    -1415181.08488224,
  
    -95475.824696437, 
    -1582706.494101,
  
    -38639.5004069032, 
    -1876739.65674409,
  
    -130158.227325917, 
    -2861634.30819273,
  
    149174.439558676, 
    -1064640.88861117,
  
    -61443.992200203, 
    -2750542.93939386,
  
    229662.746114291, 
    -2227958.50399161,
  
    121637.269316345, 
    -2824685.7916016,
  
    -242670.738696097, 
    -966680.481587737,
  
    99103.9176387681, 
    -2450775.25920432,
  
    -131530.022807945, 
    -1016997.31934229,
  
    221840.311597415, 
    -2692465.40490015,
  
    -351066.467255495, 
    -1356249.21737432,
  
    -272032.866792847, 
    -955214.885084514,
  
    243757.459174528, 
    -1180005.65926332,
  
    15951.7075890699, 
    -3040205.9110003,
  
    100030.733887794, 
    -1690121.08198604,
  
    89035.1326388729, 
    -2016305.36502083,
  
    216125.16010092, 
    -931590.38428369,
  
    48567.9136862537, 
    -2627631.50766255,
  
    225549.993284714, 
    -1826706.89785795,
  
    535282.265898878, 
    -1393361.69314196,
  
    510995.406377622, 
    -1255345.96593866,
  
    -177540.011535108, 
    -1506414.46605613,
  
    -160002.413692843, 
    -1873909.41222294,
  
    336008.371425454, 
    -2544103.00170443,
  
    -135533.275530165, 
    -3137035.16307847,
  
    -26804.7845448943, 
    -1964219.6393846,
  
    426953.18055226, 
    -1153723.16401544,
  
    684397.842787926, 
    -2196561.44783732,
  
    430088.751295958, 
    -2290747.78802541,
  
    -170892.308950487, 
    -2481770.60288364,
  
    279966.428447959, 
    -1406496.59645443,
  
    -150160.726781471, 
    -975855.895829061,
  
    -460975.991451729, 
    -1167483.4512682,
  
    459124.497814936, 
    -1116693.81318745,
  
    116625.692090824, 
    -1514250.85599311,
  
    186679.138145047, 
    -1814563.42346507,
  
    464822.469124365, 
    -1034117.17151696,
  
    109517.073734768, 
    -916970.115206676,
  
    153517.249208829, 
    -2727713.32454232,
  
    -94557.4750632621, 
    -2488013.37476937,
  
    -489639.039487239, 
    -1330861.71225432,
  
    -116864.610037569, 
    -2322818.6257473,
  
    -215120.827671591, 
    -1220790.21573909,
  
    31310.214952979, 
    -3166992.13145898,
  
    -299910.519885901, 
    -1156365.48699644,
  
    281697.632354385, 
    -1674867.47061952,
  
    422058.752224515, 
    -1322337.58468433,
  
    -145929.943849026, 
    -3102017.28619799,
  
    -119780.413449006, 
    -1672381.58556516,
  
    -121855.474890598, 
    -2068709.92801959,
  
    324730.870012546, 
    -994477.851014973,
  
    645636.722497777, 
    -2132243.77566987,
  
    23146.4486276115, 
    -1898497.34912606,
  
    174410.398310866, 
    -2799924.11967817,
  
    721902.951491267, 
    -2090874.21312104,
  
    -323180.798016995, 
    -1142063.84777306,
  
    533476.033096588, 
    -1505401.29886225,
  
    180051.596089469, 
    -1942855.34212067,
  
    65974.8478016777, 
    -2997658.22493864,
  
    302169.569576639, 
    -2261182.03629456,
  
    -59656.8231703026, 
    -2584086.79214144,
  
    66599.3119183167, 
    -1450224.88628356,
  
    -222947.814440486, 
    -2899606.16200512,
  
    -56362.1213794579, 
    -2618402.08608265,
  
    335024.622428283, 
    -1443762.73171393,
  
    411997.779152093, 
    -1752387.18992747,
  
    439376.277056687, 
    -2483173.45300319,
  
    -2674.69430312006, 
    -2658531.46092086,
  
    138565.862211675, 
    -961994.641789492,
  
    343115.760510479, 
    -1897522.21362421,
  
    307624.373602522, 
    -2240574.0416366,
  
    -470571.80395052, 
    -1180797.54127271,
  
    31365.7802942913, 
    -3146726.70992275,
  
    173394.651493967, 
    -2482209.96574568,
  
    -298711.632535678, 
    -1424583.11213621,
  
    -107019.665977631, 
    -3059502.69491349,
  
    -320431.680871945, 
    -1161476.5783042,
  
    563174.370379126, 
    -1421444.67124808,
  
    19715.1290899227, 
    -1666693.46517295,
  
    -315187.588691488, 
    -1687355.08829799,
  
    -49394.862309238, 
    -2062143.39756326,
  
    -172896.959063654, 
    -1968031.92612435,
  
    753675.611413202, 
    -2086631.98320969,
  
    40860.4389503478, 
    -2746585.94475135,
  
    -39665.0659673782, 
    -2469334.57157701,
  
    -276192.340920331, 
    -1397317.08502621,
  
    -383182.806491224, 
    -1366109.26558835,
  
    562740.449292942, 
    -1623445.67110925,
  
    386907.974010729, 
    -1921491.04265913,
  
    -19991.865850755, 
    -2870034.39136621,
  
    157357.013521745, 
    -1096491.7576947,
  
    90675.6951079902, 
    -2224875.33427813,
  
    -334006.951223056, 
    -1469678.05265437,
  
    143548.321661916, 
    -2651752.97647854,
  
    474430.409652213, 
    -1310553.17039836,
  
    -146767.804869507, 
    -1493953.17365819,
  
    541430.127473888, 
    -2207302.87760079,
  
    142297.16389382, 
    -2705369.61267378,
  
    399875.565574078, 
    -1409461.82464537,
  
    380902.455908725, 
    -1753709.7801278,
  
    353665.656579484, 
    -2537572.74646545,
  
    -190911.953479715, 
    -2592752.91982704,
  
    121080.722732177, 
    -2954164.94841913,
  
    140581.215682837, 
    -1928728.82752396,
  
    357056.0760641, 
    -1045262.82314881,
  
    103552.450923356, 
    -2179939.58078796,
  
    557399.894228357, 
    -2033999.30523575,
  
    549893.806267858, 
    -1564879.91033693,
  
    -38252.3195213462, 
    -3047012.72649523,
  
    -363841.611472135, 
    -1383558.83064491,
  
    -333437.004591125, 
    -1096923.28104516,
  
    -219501.718501582, 
    -1659229.76267795,
  
    -344666.850726992, 
    -1550677.85984466,
  
    -15115.3284717333, 
    -2968404.33752023,
  
    -268916.947219088, 
    -1882828.34049031,
  
    172501.815404436, 
    -2023532.59895626,
  
    -4567.75609768621, 
    -2721331.72686268,
  
    -235108.074100717, 
    -999670.202725039,
  
    -104655.850781123, 
    -2142748.63008765,
  
    -319339.972021325, 
    -1306186.91336532,
  
    179612.805923097, 
    -2534699.84344276,
  
    -177799.442655003, 
    -1197702.87334124,
  
    -84520.9294877598, 
    -2822313.38106669,
  
    -353980.478481945, 
    -1057017.08638655,
  
    -201532.869868273, 
    -2937980.39934289,
  
    164853.897005949, 
    -2847086.74245182,
  
    -37729.964868737, 
    -954279.883011362,
  
    -127573.420849884, 
    -2187408.97512889,
  
    463995.963895444, 
    -1719494.29375796,
  
    420491.103191471, 
    -1933941.3102671,
  
    -259269.848601366, 
    -1911241.78981525,
  
    522438.86900154, 
    -1790105.59264934,
  
    -463001.860836527, 
    -1389821.79223611,
  
    175369.951518022, 
    -1447158.09405352,
  
    167097.715886693, 
    -1801221.37129765,
  
    480874.428298894, 
    -2361177.02004565,
  
    576018.731635512, 
    -1997990.33618847,
  
    -77718.0135108529, 
    -2864550.09622332,
  
    -61953.3291447583, 
    -1959935.44142311,
  
    662502.233610874, 
    -2195962.65695124,
  
    -106171.55210755, 
    -2117625.75512854,
  
    34770.0908265139, 
    -2503424.16302243,
  
    54623.8187193043, 
    -2284260.72372157,
  
    222722.142767572, 
    -2711214.9991814,
  
    161983.451672396, 
    -2646290.40112734,
  
    493341.965513533, 
    -1451137.82291595,
  
    -522057.115234197, 
    -1375031.55381966,
  
    -443519.059450368, 
    -1183863.26701935,
  
    -225264.863769301, 
    -1624595.82822516,
  
    -177297.127013672, 
    -1915001.95578558,
  
    -4619.02828044172, 
    -2929790.14400122,
  
    281388.064409667, 
    -1171374.61186389,
  
    402498.702743342, 
    -1983512.33836284,
  
    -201879.82414904, 
    -2765457.70229167,
  
    103859.991426369, 
    -2195894.36752694,
  
    501048.460989018, 
    -2180005.87659404,
  
    -9632.2801727775, 
    -2809785.25449965,
  
    -280408.766549205, 
    -1097554.65485955,
  
    218707.953048534, 
    -2521638.03700041,
  
    -75996.8560680936, 
    -991171.277599072,
  
    136859.775665561, 
    -2829148.17069619,
  
    3883.70644769482, 
    -2982692.64746708,
  
    131523.151099565, 
    -1090412.78492124,
  
    172563.563423802, 
    -2857707.17555662,
  
    238684.154012482, 
    -1701310.87691597,
  
    216901.566871616, 
    -1984531.61743134,
  
    472111.799594868, 
    -1021947.58640033,
  
    -83264.9796912392, 
    -2589070.54449275,
  
    352942.304451602, 
    -1781522.15811711,
  
    137315.80808165, 
    -2925957.41364452,
  
    -44594.3662112596, 
    -1484091.84051035,
  
    -38223.95731203, 
    -1846847.85988319,
  
    97363.9492208435, 
    -905451.897874633,
  
    -154101.017211028, 
    -1977366.89964672,
  
    748332.845381163, 
    -2069162.0748672,
  
    -231138.706310116, 
    -2696469.76634339,
  
    294233.348727149, 
    -2288400.55767043,
  
    -438743.711023534, 
    -1406486.56969194,
  
    -37705.3429665933, 
    -2547596.6398432,
  
    529624.697320402, 
    -1288498.85514559,
  
    411269.269886106, 
    -1379586.8807302,
  
    -254734.03660058, 
    -1023953.90799238,
  
    555488.949671324, 
    -1437134.84814152,
  
    -14357.6753726981, 
    -1556525.65935273,
  
    48021.5139931468, 
    -1852825.72224912,
  
    -210836.279306654, 
    -2835383.25893493,
  
    66540.9243340568, 
    -997932.311546291,
  
    528357.020533119, 
    -2202262.44794611,
  
    23158.2443250424, 
    -2741557.8949041,
  
    -429871.250502419, 
    -1387820.61210837,
  
    19291.0513259064, 
    -2403487.87940676,
  
    -163680.332032809, 
    -1095379.2021543,
  
    282058.255567674, 
    -2633669.19172429,
  
    -331391.102783334, 
    -1279370.86048093,
  
    57160.9997228047, 
    -877590.048267068,
  
    455357.078964815, 
    -1680285.74576551,
  
    312334.880373347, 
    -1234748.70780046,
  
    -499093.417945005, 
    -1376938.49220099,
  
    -64333.5950734135, 
    -3061832.20099317,
  
    15437.0720202732, 
    -1683294.08892171,
  
    7923.36223158086, 
    -2036460.96618458,
  
    127616.718815038, 
    -2650753.18629068,
  
    146363.342555334, 
    -1854793.58747761,
  
    453940.587311199, 
    -1046369.57925839,
  
    -260631.038053551, 
    -1520366.1065219,
  
    -235343.441104152, 
    -1890651.66068975,
  
    32917.4181135645, 
    -3211310.12550999,
  
    -236591.504463194, 
    -1951440.74080498,
  
    52755.3609682361, 
    -1956002.60264126,
  
    -283002.605526636, 
    -1130319.65733845,
  
    -189991.645684511, 
    -2540686.01783175,
  
    479287.4601418, 
    -1228072.22546968,
  
    197902.153356426, 
    -1423315.17055895,
  
    -187443.759852245, 
    -2561018.1798328,
  
    200625.282113558, 
    -1487140.03804841,
  
    273340.154742136, 
    -1790649.48625678,
  
    28111.641956729, 
    -3180686.03365139,
  
    113163.619572097, 
    -2699010.56460188,
  
    5700.86026704819, 
    -928750.712729086,
  
    467752.403202834, 
    -1878318.14451573,
  
    -292518.823355865, 
    -1823539.88215218,
  
    432518.913265387, 
    -2277683.08173575,
  
    -5823.85040592671, 
    -2506636.45174275,
  
    -488004.160783134, 
    -1393820.19899182,
  
    107100.337051202, 
    -3067037.31788015,
  
    286163.726287137, 
    -2545108.80831402,
  
    -247271.136896676, 
    -1299172.09855141,
  
    18538.6623788179, 
    -3024709.44312161,
  
    -280235.152958735, 
    -1079487.1298451,
  
    -88915.5342549744, 
    -3124928.8501673,
  
    178069.550380208, 
    -1671634.21386485,
  
    482478.07864096, 
    -1186392.02184035,
  
    -68412.4738446522, 
    -3126951.96898995,
  
    -204291.340914418, 
    -1665561.27117745,
  
    -185903.647647414, 
    -2085896.40432297,
  
    475883.242875108, 
    -1117617.24613252,
  
    -53291.1604491037, 
    -1925608.98304844,
  
    582238.542079135, 
    -1476624.3736558,
  
    -78588.861165492, 
    -3173734.56406418,
  
    -187370.01876982, 
    -2425304.71099076,
  
    -346745.258480762, 
    -1230052.72542433,
  
    556126.820007151, 
    -1578903.30493409,
  
    259611.741344572, 
    -1934638.30292207,
  
    -157209.260767633, 
    -2832722.72174471,
  
    283025.480757015, 
    -1188099.86321062,
  
    -189818.609293393, 
    -3064327.78964408,
  
    221631.025452359, 
    -2247356.1551128,
  
    -314576.72452497, 
    -1340398.66398731,
  
    20006.9906947754, 
    -2610614.39962636,
  
    -15464.9634312799, 
    -1467043.45793328,
  
    609244.59162177, 
    -2168291.82133341,
  
    -218865.11255411, 
    -938792.970591383,
  
    22425.5237514667, 
    -2652893.13190655,
  
    419024.209995973, 
    -1416651.91402747,
  
    498658.79329415, 
    -1728473.25297709,
  
    386932.06444141, 
    -2543554.93929231,
  
    -75073.6398616733, 
    -2633232.02105505,
  
    226186.499448872, 
    -979427.677292597,
  
    265217.858375247, 
    -1909524.75841581,
  
    410970.123186787, 
    -1171072.54617779,
  
    -577795.736524305, 
    -1166161.79465611,
  
    -330861.941760796, 
    -1502964.99494819,
  
    -161341.973217094, 
    -3087096.90889422,
  
    -337607.789077141, 
    -1249348.37557623,
  
    -436488.725173364, 
    -1232346.70031309,
  
    -74676.4432355161, 
    -1663748.39384553,
  
    -221193.659825275, 
    -2969955.06576243,
  
    436569.482820311, 
    -2542519.02382926,
  
    -296926.006455698, 
    -1764502.29193373,
  
    35923.128139239, 
    -2047297.77055082,
  
    136579.119320095, 
    -2723542.70814118,
  
    -255388.463605774, 
    -1006894.84325586,
  
    -42560.2608181441, 
    -2759428.01309936,
  
    -343297.636310725, 
    -1434575.99412129,
  
    47793.5507981937, 
    -2495405.4023923,
  
    -238675.827765755, 
    -1321205.60367475,
  
    466468.119523793, 
    -1913274.0059153,
  
    63181.0065568843, 
    -2892650.4645162,
  
    80461.9266217462, 
    -1040437.81348702,
  
    6733.72697485245, 
    -2210465.19542833,
  
    496297.316790073, 
    -2344537.50645164,
  
    218868.798217954, 
    -2676834.2789085,
  
    -228832.080219209, 
    -1510771.74530805,
  
    -212924.52044251, 
    -2018186.6606743,
  
    -205630.667250607, 
    -2320840.88306978,
  
    313527.253707907, 
    -1423960.39062743,
  
    297338.755659877, 
    -1772279.26702191,
  
    418060.863452527, 
    -2485573.20411556,
  
    -219344.958848606, 
    -2676368.11498468,
  
    50752.6382077565, 
    -2909423.78252494,
  
    62683.3135476012, 
    -1940731.37231535,
  
    22889.3714134532, 
    -2155972.72396004,
  
    -105266.404773338, 
    -2281498.23233578,
  
    522089.548287104, 
    -1490678.3761419,
  
    36894.8679340138, 
    -3022541.02552768,
  
    -379462.930822584, 
    -1463476.43667006,
  
    -349115.789412008, 
    -1076578.35354017,
  
    -331656.107990578, 
    -1603857.79395132,
  
    413601.6892613, 
    -1278108.33511693,
  
    260962.158338365, 
    -2008140.19219898,
  
    -101058.997424831, 
    -2719820.25023778,
  
    -24457.449474923, 
    -2163189.29904944,
  
    527032.408176687, 
    -2046346.05272558,
  
    -146598.11981924, 
    -2794238.12646035,
  
    -304366.430838676, 
    -1225943.73561558,
  
    -138644.601759177, 
    -1118267.64326524,
  
    2428.1885330317, 
    -2824997.80226872,
  
    -121875.035294577, 
    -2955319.21926626,
  
    41737.5073834622, 
    -3098527.97733606,
  
    18275.7030983384, 
    -1000011.15664478,
  
    377337.576592179, 
    -1712500.67158778,
  
    342187.435783898, 
    -1953399.11914465,
  
    514327.516323829, 
    -2200772.03763627,
  
    483381.257333341, 
    -1735256.80543158,
  
    -457129.331100759, 
    -1293329.36478731,
  
    89021.6369388325, 
    -1461656.65783883,
  
    87169.4528580752, 
    -1818982.99334812,
  
    463664.226276504, 
    -2319237.15748457,
  
    528610.617618254, 
    -1819091.18299486,
  
    -139851.231279923, 
    -1971937.98621421,
  
    635292.000202326, 
    -2116746.08954925,
  
    -61010.2947107252, 
    -2479127.61188306,
  
    149732.544601748, 
    -2285903.95605727,
  
    87438.2353923384, 
    -2609447.33371722,
  
    505997.423217344, 
    -1551012.26393636,
  
    686467.819140595, 
    -2107805.99050676,
  
    568615.715773232, 
    -1438093.67120789,
  
    411843.564209204, 
    -2400482.76254416,
  
    -144146.714187482, 
    -1598414.99593197,
  
    -90636.1104167144, 
    -1891088.01857782,
  
    -82430.7876521992, 
    -2887545.76499714,
  
    198754.549184592, 
    -1104666.03479862,
  
    490959.042964153, 
    -1968119.92940818,
  
    -113065.448901098, 
    -2756025.31249903,
  
    182845.565378962, 
    -2216025.91518162,
  
    485497.357591565, 
    -2259999.79561768,
  
    73325.0098140666, 
    -2819201.82012856,
  
    541074.287147753, 
    -1643460.16561932,
  
    145047.959267923, 
    -2477996.09864319,
  
    -112239.836136249, 
    -969968.191025003,
  
    -468095.828939022, 
    -1349985.74455313,
  
    -362871.688135768, 
    -1402376.23422336,
  
    185878.01643537, 
    -2860118.07284595,
  
    202302.805987241, 
    -1146913.8044678,
  
    64122.8886956854, 
    -3027230.13705588,
  
    152025.766709176, 
    -1694317.25474563,
  
    137702.196898897, 
    -2004212.00460708,
  
    -176.916981613265, 
    -2613373.70300329,
  
    273110.471838109, 
    -1809837.68582849,
  
    592174.066852627, 
    -2012170.4441754,
  
    -127685.395184664, 
    -1498043.48123408,
  
    -114797.798667443, 
    -1863864.06378861,
  
    360310.770464185, 
    -2501294.31941961,
  
    -84418.5766721066, 
    -3151867.32905876,
  
    -74540.8716979416, 
    -1969149.86290356,
  
    679061.024087602, 
    -2146041.38544244,
  
    380233.298721648, 
    -2289886.4142439,
  
    -456505.860946616, 
    -1314036.64023482,
  
    -120061.416216322, 
    -2506893.15196315,
  
    536012.936468282, 
    -1918860.67993245,
  
    329204.994794538, 
    -1396405.45483458,
  
    -194511.681029294, 
    -997419.979365965,
  
    431611.220254268, 
    -1070984.14522923,
  
    66760.4739510061, 
    -1530344.82460448,
  
    134682.528135191, 
    -1828911.785299,
  
    568989.286332207, 
    -2104021.45121347,
  
    105449.279267653, 
    -2732818.30672415,
  
    -149302.994639994, 
    -2476523.59176892,
  
    -479229.453072214, 
    -1376124.78100409,
  
    -64353.7214826615, 
    -2353930.17896493,
  
    -195830.641257774, 
    -1173761.08496649,
  
    -311715.738311165, 
    -1202492.5035875,
  
    67499.9843597369, 
    -888647.763259333,
  
    345676.317316436, 
    -1676863.64302065,
  
    380912.301572314, 
    -1289491.75633763,
  
    -144618.895280561, 
    -3083458.49072737,
  
    -69073.855445138, 
    -1676473.77453398,
  
    -73188.4106306736, 
    -2056616.56760615,
  
    283322.44150364, 
    -972448.739132458,
  
    203898.911262964, 
    -2673065.63496213,
  
    69352.7849001497, 
    -1882108.43963868,
  
    505430.775759662, 
    -1227372.72416193,
  
    735761.423718259, 
    -2127126.77904744,
  
    -308646.279317192, 
    -1087792.45634986,
  
    519564.289902865, 
    -1460257.56094511,
  
    132315.50867837, 
    -1947785.56318477,
  
    17896.6595279135, 
    -2989439.98706433,
  
    -295146.497826779, 
    -1211119.27531999,
  
    -107882.894280288, 
    -2568027.77747774,
  
    115837.878006859, 
    -1440133.74220854,
  
    -104263.978847406, 
    -2597431.9803062,
  
    284624.869681247, 
    -1460029.22036182,
  
    360001.169142234, 
    -1766735.55176149,
  
    471686.122202003, 
    -2445973.61141582,
  
    40764.6740139173, 
    -2673711.12473689,
  
    82754.9632145945, 
    -950890.483832592,
  
    389854.501067635, 
    -1890320.68930746,
  
    79494.7472283913, 
    -2524542.7947415,
  
    -485946.553823636, 
    -1225705.99936328,
  
    216934.07150717, 
    -2506494.80749476,
  
    -279421.446121801, 
    -1377553.98136369,
  
    -59935.2945885575, 
    -3046455.22660588,
  
    -309703.632005159, 
    -1106592.61441009,
  
    516055.167211137, 
    -1405006.28457336,
  
    78011.3789392012, 
    -1668512.34182374,
  
    491087.404540822, 
    -1276487.41007898,
  
    204755.20875164, 
    -2876824.88740284,
  
    -556470.260614352, 
    -1370197.96555271,
  
    -288802.268379832, 
    -1658740.95678975,
  
    -100585.65745709, 
    -2071050.77485585,
  
    573369.50858151, 
    -2258685.49938827,
  
    -128044.784712238, 
    -1952123.32124344,
  
    717894.50216551, 
    -2071799.58882377,
  
    90155.625229135, 
    -2738997.27418936,
  
    -93799.3934380694, 
    -2453197.4904043,
  
    -298702.250440922, 
    -1442983.97251881,
  
    -369674.866429238, 
    -1315671.08593892,
  
    592670.154461078, 
    -1525741.31502685,
  
    339171.886857691, 
    -1926421.26617839,
  
    203496.210117094, 
    -1130125.68646967,
  
    141040.875057419, 
    -2233521.4181821,
  
    -326720.616825048, 
    -1421198.28196879,
  
    97590.253657075, 
    -2636449.19559518,
  
    573899.49213942, 
    -2157029.35504071,
  
    98127.7896584862, 
    -2686033.48469353,
  
    451684.555897865, 
    -1400762.68720156,
  
    -147472.585162382, 
    -2607932.58364381,
  
    307415.96743757, 
    -995589.124999897,
  
    187319.956240005, 
    -1921527.30320733,
  
    376553.415070727, 
    -1090760.33137628,
  
    151506.198409355, 
    -2194187.74157568,
  
    547376.410081281, 
    -1977663.188961,
  
    -517466.374050319, 
    -1183659.6375226,
  
    547242.47924683, 
    -1624934.15591474,
  
    -84386.7622276874, 
    -3062036.42271561,
  
    -354181.493294856, 
    -1334138.32230464,
  
    -370070.879904252, 
    -1145064.97634737,
  
    -165812.50696352, 
    -1660904.89795511,
  
    554188.82582452, 
    -1852340.43002266,
  
    -279228.228664163, 
    -1839267.67733927,
  
    121241.120784752, 
    -2032452.14082515,
  
    50129.5252209155, 
    -2722188.52637232,
  
    -192207.776293221, 
    -954082.76228376,
  
    -152774.890634471, 
    -2130484.22811625,
  
    230594.751992332, 
    -927617.064628328,
  
    -128430.644021241, 
    -2772647.19299057,
  
    -328324.09512813, 
    -1354332.81637169,
  
    -201159.314353196, 
    -1245094.12477825,
  
    -137690.777544964, 
    -2820671.84417321,
  
    149566.993170951, 
    -2897837.6715374,
  
    6591.99434337548, 
    -986589.106019025,
  
    -77208.2384453053, 
    -2196055.05877525,
  
    558191.064153599, 
    -2089830.30482909,
  
    527071.54625807, 
    -1837823.62300327,
  
    -96106.893315642, 
    -3139548.51570136,
  
    227178.939128705, 
    -1438458.95441259,
  
    215938.107707414, 
    -1790368.08261449,
  
    482060.340731736, 
    -2415459.93488958,
  
    -28654.9783897729, 
    -2881687.38867462,
  
    -15214.5885876169, 
    -1952733.91710663,
  
    776877.636676347, 
    -2042165.13634915,
  
    -57773.7053835059, 
    -2132005.86932882,
  
    -4340.01449122214, 
    -2283241.97979601,
  
    492318.155382931, 
    -1411227.11931093,
  
    345750.49598342, 
    -2507079.98266279,
  
    -273935.750805338, 
    -1640304.32979803,
  
    -229293.734568387, 
    -1929350.31736108,
  
    41469.8352491811, 
    -2954812.00965884,
  
    330968.174035843, 
    -1211399.75805151,
  
    349422.498559229, 
    -1992747.78324457,
  
    -204508.904453633, 
    -2718199.77121363,
  
    -584297.990057454, 
    -1152981.99888704,
  
    55740.9518311905, 
    -2183629.96801097,
  
    510597.667473803, 
    -2130885.3441859,
  
    -60465.0973903441, 
    -2804015.17037565,
  
    -289392.891853012, 
    -1145700.56057892,
  
    261165.680295807, 
    -2546793.31103572,
  
    -99489.7606054454, 
    -1038832.41564445,
  
    87225.1454199583, 
    -2827615.77721858,
  
    -544786.676605607, 
    -1170140.69497895,
  
    -42680.7478048064, 
    -2972557.13866891,
  
    597813.183943984, 
    -1549272.86396684,
  
    89055.3579856921, 
    -1056512.17619103,
  
    -508126.656602921, 
    -1196204.50318688,
  
    25099.7286084995, 
    -3108631.28906953,
  
    290679.186833861, 
    -1705507.04967554,
  
    263883.768634355, 
    -1972856.93047711,
  
    485102.839915789, 
    -2276669.90711307,
  
    401856.911071735, 
    -1764172.65000392,
  
    5260.25039718336, 
    -1475720.85814337,
  
    8798.57150175426, 
    -1836398.53493256,
  
    424438.87799115, 
    -2388332.62733591,
  
    47116.2919684583, 
    -901822.810990911,
  
    -201837.104364037, 
    -1982297.12316557,
  
    649731.311520132, 
    -2183693.53106924,
  
    770874.458401043, 
    -2065765.13074191,
  
    -163216.906014823, 
    -2453200.92306945,
  
    241088.311402911, 
    -2287482.34894549,
  
    -458952.34958249, 
    -1371433.34214449,
  
    10146.3785052074, 
    -2571246.77322962,
  
    519763.427185032, 
    -1659650.91922193,
  
    460507.836232716, 
    -1369495.73911043,
  
    -213646.336468913, 
    -995735.281612866,
  
    454037.814975829, 
    -2332430.39099857,
  
    -63028.5648637237, 
    -1572234.1611837,
  
    -3975.09627472297, 
    -1867174.08162792,
  
    116121.033959799, 
    -1037957.45773357,
  
    -27029.6879049346, 
    -2746888.02235362,
  
    260874.198129103, 
    -2235913.56173354,
  
    153845.443308196, 
    -2828341.7741342,
  
    -209606.899711692, 
    -947956.034476428,
  
    67745.4346670889, 
    -2432196.04271563,
  
    -144390.145361047, 
    -1048350.07383687,
  
    197655.146467449, 
    -2713695.13803033,
  
    -343196.321466633, 
    -1325497.87461698,
  
    -245238.08870974, 
    -928544.948781589,
  
    271188.427266244, 
    -1201902.87971179,
  
    -16162.413966963, 
    -3048856.42704913,
  
    66143.6300241429, 
    -1687386.27789054,
  
    56590.4240365516, 
    -2024367.60602897,
  
    183252.694890989, 
    -917508.821930947,
  
    80498.0258591007, 
    -2636971.02700354,
  
    193843.006764111, 
    -1837953.03929692,
  
    -210776.421703081, 
    -1511995.12169982,
  
    -190138.826078781, 
    -1880606.3122555,
  
    5019.27355714238, 
    -1960932.82370527,
  
    415229.776544494, 
    -1114222.71360469,
  
    701991.441444211, 
    -2155427.31832781,
  
    462932.493814565, 
    -2291315.24224172,
  
    479536.86502495, 
    -1289323.51359519,
  
    247140.719444962, 
    -1413224.02648402,
  
    -120593.425586307, 
    -961479.840309844,
  
    -462423.918284037, 
    -1204289.20231404,
  
    150225.529624543, 
    -1503406.5291514,
  
    221343.544732275, 
    -1804997.84809076,
  
    156602.987888884, 
    -2714190.22841741,
  
    69359.6764359714, 
    -921526.997190748,
  
    514491.143501925, 
    -1871116.61774387,
  
    -276295.439420766, 
    -1867825.08957888,
  
    -58711.2397717033, 
    -2495536.64653416,
  
    -152768.857672196, 
    -2301546.1450256,
  
    -227980.950482821, 
    -1252142.96777879,
  
    65623.0362231856, 
    -3011661.97455537,
  
    -136568.090885801, 
    -3112208.99968847,
  
    239836.449354968, 
    -1673561.37784542,
  
    449489.72277139, 
    -1344234.80487475,
  
    -115126.873316778, 
    -3111925.56587822,
  
    -153584.782910548, 
    -1669653.46014626,
  
    -154300.183492841, 
    -2076772.1690275,
  
    661872.213828967, 
    -2164891.13434007,
  
    -7657.77546806107, 
    -1909423.28960262,
  
    -131812.057639521, 
    -3172676.93711352,
  
    693416.352171633, 
    -2074974.85971071,
  
    -332648.923655976, 
    -1177417.49394034,
  
    542536.348791235, 
    -1534802.10069682,
  
    211875.654191512, 
    -1939568.52644124,
  
    -147.106408555984, 
    -914263.066294739,
  
    269954.151332728, 
    -2255651.68289149,
  
    -307290.390126913, 
    -1291918.89330158,
  
    418430.833046256, 
    -1088574.24209507,
  
    33773.6026572783, 
    -1456952.31385821,
  
    611620.960047312, 
    -2230600.99177925,
  
    -264029.558331832, 
    -974678.809900154,
  
    -24427.548915877, 
    -2632382.15651414,
  
    368624.457506964, 
    -1432918.40513034,
  
    446662.183284295, 
    -1742821.61481114,
  
    418208.747201073, 
    -2507544.62482176,
  
    -31634.2715445064, 
    -2648411.68487138,
  
    174448.695406387, 
    -969133.903953496,
  
    311956.598674377, 
    -1902323.23164407,
  
    432923.749345283, 
    -1222301.85768557,
  
    276400.738072949, 
    -2231296.78167615,
  
    161871.13184958, 
    -2541831.63777391,
  
    68709.9927541886, 
    -3131154.62168109,
  
    143702.853618149, 
    -2465648.86734724,
  
    -311571.755346933, 
    -1455935.86417582,
  
    -138409.24935864, 
    -3068201.00737647,
  
    -327368.324066924, 
    -1196963.97406707,
  
    547381.284817534, 
    -1409153.96753668,
  
    -18628.0466742703, 
    -1665497.13577047,
  
    647716.940753563, 
    -2259923.42271808,
  
    -307782.155534829, 
    -1718639.80301553,
  
    -15267.6670086509, 
    -2056205.14784354,
  
    35771.562611775, 
    -879647.971773937,
  
    726264.548897076, 
    -2061743.9681841,
  
    7867.13318120767, 
    -2751665.04794342,
  
    -352281.759159445, 
    -1482721.8995825,
  
    -4231.1005024604, 
    -2479897.20187889,
  
    -261185.737028298, 
    -1366872.49362247,
  
    -391996.107314506, 
    -1399017.82422721,
  
    418732.032112747, 
    -1918204.2269796,
  
    13351.0558787094, 
    -2879100.87924261,
  
    126597.548134528, 
    -1074069.13696076,
  
    57098.9093793687, 
    -2219111.27907443,
  
    511061.84311675, 
    -2236019.02287511,
  
    -203478.567973032, 
    -2360396.63634417,
  
    365336.24131861, 
    -1415261.25098658,
  
    347130.320221968, 
    -1761214.60982241,
  
    379423.739044098, 
    -2516772.93154122,
  
    -210587.522627861, 
    -2620713.11416701,
  
    98397.2095359099, 
    -2926065.61769796,
  
    109422.053846731, 
    -1933529.84554374,
  
    344613.365077632, 
    -1016227.45893302,
  
    71287.2181374006, 
    -2170352.83816004,
  
    -8193.44355722678, 
    -3037224.04600507,
  
    -370163.537036304, 
    -1415901.36556858,
  
    18609.5218539824, 
    -2974052.95391362,
  
    207885.95169921, 
    -2017375.63733859,
  
    -42374.3549349489, 
    -2720739.50994617,
  
    -72576.489328231, 
    -2150924.89707818,
  
    537222.833568287, 
    -1993927.12590471,
  
    -199301.029766235, 
    -2788255.7652078,
  
    -313350.556142487, 
    -1274089.64133502,
  
    -162137.506296658, 
    -1165928.78131082,
  
    -49486.6054054204, 
    -2823395.01134193,
  
    125727.640385854, 
    -3068520.48614159,
  
    -169669.73544456, 
    -2944915.92824271,
  
    -24192.0900153474, 
    -966110.547914783,
  
    -161150.206578573, 
    -2181644.91992492,
  
    429332.60941354, 
    -1716696.84434729,
  
    389169.635349647, 
    -1941724.43490336,
  
    532564.373164158, 
    -2153410.0518034,
  
    140830.624549516, 
    -1452957.51819783,
  
    134537.457299927, 
    -1808456.89846506,
  
    480114.397978417, 
    -2326387.99518263,
  
    -258354.169630946, 
    -2894455.2079677,
  
    -93112.4909808396, 
    -1964736.45944278,
  
    -138436.784635577, 
    -2108039.01495535,
  
    92869.5401667929, 
    -2284921.50930036,
  
    132567.340167094, 
    -2631751.8454586,
  
    498276.41965547, 
    -1490079.58930433,
  
    726601.242191588, 
    -2139808.26086723,
  
    -453669.406553268, 
    -1224475.29753398,
  
    386790.003222976, 
    -2440890.02381367,
  
    -192817.603936571, 
    -1614123.49530789,
  
    -142632.720426504, 
    -1905436.38041149,
  
    -35344.9388509591, 
    -2913108.90121966,
  
    248334.658810609, 
    -1144691.18098615,
  
    437882.838780066, 
    -1977355.37428999,
  
    -166281.06100664, 
    -2761676.99296594,
  
    135939.35313719, 
    -2204070.6369722,
  
    494711.846303587, 
    -2212601.03440527,
  
    23551.6050585383, 
    -2813551.99135211,
  
    -274419.350412335, 
    -1065457.38528435,
  
    189810.739269454, 
    -2504517.06835298,
  
    -60334.919709888, 
    -959397.185568877,
  
    -374676.906819032, 
    -1448503.24835927,
  
    34926.6765096301, 
    -2989449.65079139,
  
    611453.949578776, 
    -1530576.40185564,
  
    159835.012615212, 
    -1113013.19328245,
  
    75912.0722517631, 
    -3044308.66871112,
  
    204020.799530558, 
    -1698513.42750523,
  
    185580.101484819, 
    -1992314.74180944,
  
    -50029.7560287722, 
    -2598791.80854286,
  
    320670.95284653, 
    -1792968.47354096,
  
    -77830.7788342338, 
    -1489672.49641204,
  
    -69572.3123095737, 
    -1853814.07677495,
  
    384613.166789916, 
    -2458485.63493733,
  
    132090.20765921, 
    -907959.969734828,
  
    -122276.959109011, 
    -1974080.08396746,
  
    462123.393091618, 
    -1272224.52015781,
  
    329027.947070252, 
    -2289001.71885977,
  
    -445299.340282971, 
    -1372365.27539418,
  
    -70360.3332881793, 
    -2531457.30946623,
  
    378443.558428066, 
    -1386314.31101777,
  
    -238862.633080191, 
    -1018984.06018987,
  
    18089.584460001, 
    -1546053.32643544,
  
    82685.9205803654, 
    -1843260.14687487,
  
    -213100.914931089, 
    -2869252.67784782,
  
    33487.5187352929, 
    -971248.880668823,
  
    544038.256491931, 
    -2164348.2408852,
  
    56388.065480884, 
    -2738028.77518488,
  
    338902.828424026, 
    -2255801.20854315,
  
    -13624.313001487, 
    -2383986.24466511,
  
    -176540.454585954, 
    -1126731.95664896,
  
    -323520.956994467, 
    -1248619.51772356,
  
    410715.770800476, 
    -1678892.91164721,
  
    339765.848207092, 
    -1256645.92579392,
  
    -96447.7141743019, 
    -3070482.71678372,
  
    -18367.2974412693, 
    -1680565.9635028,
  
    -24521.3488257436, 
    -2044523.20745066,
  
    240663.105400185, 
    -949754.147892069,
  
    158364.6492911, 
    -2659746.9189009,
  
    115559.118459641, 
    -1865719.52795426,
  
    185508.333111106, 
    -2789477.15406616,
  
    -293867.44822154, 
    -1525946.76216559,
  
    539694.88430212, 
    -2279127.15260481,
  
    505573.156805672, 
    -1414856.21025764,
  
    84579.4190702786, 
    -1952715.78696189,
  
    -32778.5645469175, 
    -2980777.82763943,
  
    398815.821337088, 
    -2277773.09185141,
  
    -287860.163428703, 
    -1162639.50463427,
  
    -157148.145071194, 
    -2551622.72218122,
  
    165076.444095397, 
    -1430042.59813355,
  
    -561159.013451082, 
    -1170649.08027235,
  
    -154130.028778506, 
    -2575602.00690696,
  
    234225.117192241, 
    -1476295.71146477,
  
    308004.559132373, 
    -1781083.9135955,
  
    468728.303034808, 
    -2481217.65331994,
  
    84204.0398758416, 
    -2688890.78881077,
  
    24350.6839744225, 
    -939270.345661191,
  
    436593.241366747, 
    -1883119.16253564,
  
    -303334.411741567, 
    -1794016.41126658,
  
    -484315.421846933, 
    -1189207.21369018,
  
    89621.0495088371, 
    -3052113.70182861,
  
    258866.611057865, 
    -2529883.38577866,
  
    -260131.259707926, 
    -1330524.85059111,
  
    -56024.6991774107, 
    -3133708.37019158,
  
    137706.858369221, 
    -1670374.87665793,
  
    -238095.712830986, 
    -1662833.14601659,
  
    -83192.610102759, 
    -1936214.71881747,
  
    -149352.035774176, 
    -2436637.61850154,
  
    -321212.157506484, 
    -1488650.85975329,
  
    -356016.720522262, 
    -1264672.03726354,
  
    573462.248574521, 
    -1566458.75025805,
  
    291435.799446609, 
    -1931351.4872426,
  
    251054.563228529, 
    -1164794.13424778,
  
    -198958.875013362, 
    -3028568.24942242,
  
    189415.607466419, 
    -2241825.80416464,
  
    -319434.282427017, 
    -1372718.51128314,
  
    443270.631353335, 
    -1187037.69003994,
  
    -235768.168169894, 
    -943761.493864248,
  
    53027.26890072, 
    -2666289.72766609,
  
    404689.814017598, 
    -2540643.43686458,
  
    -104033.216845105, 
    -2623112.24746041,
  
    259477.425474474, 
    -986051.2536842,
  
    234058.69653914, 
    -1914325.77643564,
  
    396931.552671158, 
    -1138313.20640337,
  
    198341.650347363, 
    -2208103.63041821,
  
    241291.988574429, 
    -2558500.18794591,
  
    557292.782927857, 
    -2016391.68724095,
  
    497193.731007477, 
    -1089010.31580185,
  
    -130559.888433584, 
    -3077072.71338924,
  
    -344308.307088149, 
    -1283627.77413015,
  
    -409071.332827257, 
    -1196316.66561019,
  
    -112012.035918182, 
    -1662583.50281707,
  
    -289797.854044798, 
    -1794615.62534312,
  
    70050.3256368384, 
    -2041359.51811796,
  
    -230116.188138118, 
    -985770.0113064,
  
    -76744.5316625564, 
    -2764690.45589312,
  
    -337308.220431912, 
    -1402478.72209106,
  
    81376.1994029996, 
    -2505416.16560071,
  
    -223669.223873739, 
    -1290761.01227097,
  
    -191700.666120822, 
    -2819004.37321662,
  
    77371.2431916357, 
    -3166912.61917329,
  
    95697.1463586788, 
    -2901492.13780898,
  
    50913.9538135879, 
    -1018898.3314818,
  
    -26843.0587538043, 
    -2204701.14022451,
  
    278987.926739393, 
    -1429759.81477168,
  
    264778.497073111, 
    -1779514.79418935,
  
    443818.94591722, 
    -2464773.38919103,
  
    563580.128460398, 
    -1982759.49192972,
  
    18989.59319662, 
    -2898329.22630309,
  
    31524.151711501, 
    -1945532.39033509,
  
    -9375.85865949305, 
    -2146385.983529,
  
    141955.972553803, 
    -2530613.94220674,
  
    -64664.1659654453, 
    -2282199.73354536,
  
    259707.600278736, 
    -2640424.4672144,
  
    -380908.11855278, 
    -1092403.04112726,
  
    321126.79169137, 
    -2546793.95846272,
  
    87558.6963235952, 
    -2979833.87557415,
  
    380548.281207073, 
    -1251424.90449719,
  
    296346.294375106, 
    -2001983.22812623,
  
    -141558.131334171, 
    -2719185.85661701,
  
    7621.91197793792, 
    -2171365.56603987,
  
    520443.128486397, 
    -2080240.89664254,
  
    -111704.475622708, 
    -2798198.93685014,
  
    -298377.014701798, 
    -1193846.4660403,
  
    -122982.665142848, 
    -1086493.55368991,
  
    476134.678689119, 
    -1093408.50627568,
  
    -90011.9011289533, 
    -2962254.74571083,
  
    18174.9139468734, 
    -3122876.41965884,
  
    342674.219655237, 
    -1709703.2224351,
  
    310865.967942071, 
    -1961182.24378086,
  
    55114.8667475833, 
    -1467349.8733214,
  
    55821.1003155449, 
    -1825949.2099819,
  
    447974.087608179, 
    -2346875.34684664,
  
    624822.280766636, 
    -2138533.39912862,
  
    -101117.053298578, 
    -2468953.75567195,
  
    186455.663376098, 
    -2286538.43643915,
  
    56864.1556519142, 
    -2594336.46744903,
  
    511367.011520087, 
    -1593388.00650469,
  
    -171121.778867825, 
    -966529.837280267,
  
    541824.773332427, 
    -1422910.41429895,
  
    428721.265006847, 
    -2373261.81387444,
  
    -111699.454612795, 
    -1587942.66055965,
  
    -55971.7038295201, 
    -1881522.44320366,
  
    -114249.082404677, 
    -2870271.46063293,
  
    165701.143585646, 
    -1077982.60392096,
  
    526343.179000855, 
    -1961962.96533527,
  
    -78651.1443478295, 
    -2752370.39791395,
  
    280212.837927649, 
    -2614624.79841606,
  
    214057.017651849, 
    -2223980.97537866,
  
    105533.183547922, 
    -2822857.80020625,
  
    114783.16022308, 
    -2460064.86609209,
  
    -125099.961402383, 
    -1001320.94332253,
  
    -355001.542346916, 
    -1371624.89146605,
  
    187644.171578811, 
    -2803800.81682286,
  
    230041.973901167, 
    -1169057.04916811,
  
    32008.7671395898, 
    -3035880.65310486,
  
    117362.412227252, 
    -1691519.80533489,
  
    105257.488038532, 
    -2012274.24316023,
  
    32480.0071382399, 
    -2622925.81270259,
  
    241403.485317503, 
    -1821083.82726748,
  
    554650.687550601, 
    -1395409.22946801,
  
    -160921.805352627, 
    -1503624.13687776,
  
    -144934.208598367, 
    -1870560.96356317,
  
    344109.171191035, 
    -2529833.44176121,
  
    -117855.330038084, 
    -3142164.84640022,
  
    -42716.8135959112, 
    -1965863.04722426,
  
    432814.881457648, 
    -1173473.39057736,
  
    682586.389581643, 
    -2179413.64695368,
  
    -179612.387129575, 
    -2955678.81042945,
  
    413666.879907628, 
    -2290464.05968973,
  
    -153699.249355215, 
    -2490268.06459158,
  
    296379.283078476, 
    -1403132.88266715,
  
    -164944.377379063, 
    -983043.923588678,
  
    449660.737457559, 
    -1100971.02983156,
  
    99825.774680493, 
    -1519673.02051246,
  
    169346.934722417, 
    -1819346.20992471,
  
    416931.461173743, 
    -2275688.85509433,
  
    -112742.380967486, 
    -2484196.7958087,
  
    -99339.5497631029, 
    -2333201.84016161,
  
    -208690.76626598, 
    -1205113.83971924,
  
    50569.8839109908, 
    -3178164.74168817,
  
    -303845.592522299, 
    -1171741.16083014,
  
    106653.234558673, 
    -880794.10656096,
  
    302628.22127005, 
    -1675520.51603709,
  
    408343.269406108, 
    -1311388.97433108,
  
    -102878.227361706, 
    -1673745.64937311,
  
    38548.5608044673, 
    -1893034.38011528,
  
    498993.979457648, 
    -1261441.83267641,
  
    731679.315629228, 
    -2105115.27709272,
  
    -318335.960173087, 
    -1123973.383319,
  
    164139.566780414, 
    -1944498.74750536,
  
    318277.277213036, 
    -2263947.21067007,
  
    -300004.05327382, 
    -1243439.12235781,
  
    -75626.028418528, 
    -2578769.13573947,
  
    83012.1662908008, 
    -1446861.17004121,
  
    -72329.4063837539, 
    -2611412.05073785,
  
    318224.704759927, 
    -1449184.89377821,
  
    11805.0943175599, 
    -2663591.34894557,
  
    120368.555340849, 
    -958374.098026678,
  
    358695.338973504, 
    -1895121.70487231,
  
    323236.190010766, 
    -2245212.67051831,
  
    112999.431691742, 
    -2531574.63101901,
  
    188213.920894619, 
    -2490475.66204034,
  
    -292281.571388083, 
    -1408906.73366138,
  
    39147.2125450378, 
    -1667299.75902656,
  
    535665.7913843, 
    -2265749.26481537,
  
    -157946.234365864, 
    -1962729.05701238,
  
    -57562.439721948, 
    -2463999.48444282,
  
    -378776.157307094, 
    -1349654.98639793,
  
    370995.944959717, 
    -1923134.45049889,
  
    -36763.6787271381, 
    -2865473.85825606,
  
    172736.744729822, 
    -1107703.06573568,
  
    -214885.330665634, 
    -2988439.00795987,
  
    107464.089328824, 
    -2227757.36297846,
  
    -331578.174727073, 
    -1453518.12926454,
  
    551967.775306053, 
    -2190987.04604911,
  
    127660.757467386, 
    -2698962.19942724,
  
    397788.523752103, 
    -1749957.3652805,
  
    -176432.162403914, 
    -2597812.80759396,
  
    112001.186007424, 
    -2971169.7234347,
  
    156160.794145864, 
    -1926328.3187721,
  
    363518.717704754, 
    -1060343.55143443,
  
    119685.067316326, 
    -2184732.95210189,
  
    272166.169898814, 
    -2563644.28335034,
  
    -511383.741928939, 
    -1221319.4237258,
  
    -345372.527305126, 
    -1112608.11818502,
  
    67100.4830076164, 
    -865981.606053913,
  
    -31977.7547330977, 
    -2965580.03068003,
  
    155368.315827338, 
    -2026513.88865025,
  
    13919.2759789394, 
    -2721621.31463646,
  
    -120695.529181564, 
    -2138660.49510683,
  
    -163805.852677584, 
    -2778092.97500265,
  
    -322334.678991264, 
    -1322235.54679643,
  
    163532.173993166, 
    -2529906.31517039,
  
    -185630.410834181, 
    -1213589.91935645,
  
    -102038.090172399, 
    -2821772.56702754,
  
    159758.262480284, 
    -2864003.7196321,
  
    -110785.026629011, 
    -2190291.00382936,
  
    481327.642234888, 
    -1720893.01710676,
  
    436151.834657357, 
    -1930049.748207,
  
    551335.385857718, 
    -2104660.84083882,
  
    549791.401853087, 
    -1367833.47807805,
  
    523999.216853632, 
    -1806177.66824428,
  
    -67530.8795149033, 
    -3153791.98436243,
  
    192639.612418232, 
    -1444258.38101189,
  
    183377.846407589, 
    -1797603.60758492,
  
    481268.883740657, 
    -2379232.47842557,
  
    -61219.7693669451, 
    -2870312.78980868,
  
    667522.738749805, 
    -2210578.7423101,
  
    -90038.938169549, 
    -2122419.12670067,
  
    34969.2074771074, 
    -2283921.14077638,
  
    490919.821747525, 
    -1432022.72802538,
  
    -438854.525463763, 
    -1165200.24793126,
  
    362166.298930832, 
    -2480603.99961428,
  
    -241488.490972607, 
    -1629831.99688078,
  
    -194629.327981242, 
    -1919784.74198706,
  
    10743.9246787795, 
    -2938130.7668775,
  
    297914.765981699, 
    -1184716.32743178,
  
    384806.634595961, 
    -1986590.81917175,
  
    87820.3132840094, 
    -2191806.23500128,
  
    504231.528912931, 
    -2163632.36505905,
  
    -26305.5109977647, 
    -2807892.66012488,
  
    -283403.475716137, 
    -1113603.29100369,
  
    233156.562393074, 
    -2530198.52106604,
  
    -83827.8242472048, 
    -1007058.32361418,
  
    602983.818622699, 
    -1515075.34031514,
  
    45424.6666083555, 
    -3082902.24136571,
  
    256015.832351939, 
    -1702709.60026481,
  
    232562.300792529, 
    -1980640.05511327,
  
    -100109.952289847, 
    -2584143.41052908,
  
    369247.174143321, 
    -1775738.98866004,
  
    -27976.1622257834, 
    -1481301.51404505,
  
    -22549.7810407697, 
    -1843364.75156631,
  
    408748.739064824, 
    -2415970.81424252,
  
    80422.5198224754, 
    -904228.320362587,
  
    -170013.046262033, 
    -1979010.30748634,
  
    701307.069588777, 
    -2199438.3917454,
  
    276518.33619973, 
    -2288094.48727712,
  
    -21754.7682382932, 
    -2555480.01837104,
  
    427682.124516633, 
    -1376223.16694295,
  
    -30581.3052890498, 
    -1561761.82581138,
  
    30689.3105705222, 
    -1857608.50870872,
  
    83067.628360968, 
    -1011274.02685603,
  
    -424860.93909548, 
    -1404650.35138301,
  
    292085.650143884, 
    -2243868.61947542,
  
    35585.5815895851, 
    -2413142.03213132,
  
    -157250.270627226, 
    -1079702.82613449,
  
    -335326.175677769, 
    -1294746.53185962,
  
    477786.106539264, 
    -1680985.54480386,
  
    298619.395099953, 
    -1223800.09770524,
  
    -497641.114433359, 
    -1361989.15827336,
  
    -48276.5330679247, 
    -3057506.94283983,
  
    32339.2581075742, 
    -1684658.15272966,
  
    24145.7151762044, 
    -2032429.84458204,
  
    111959.899971151, 
    -2646173.58678304,
  
    162136.020243511, 
    -1849199.18073587,
  
    -316402.742247711, 
    -1766341.76024797,
  
    -244012.831871062, 
    -1517575.77734352,
  
    -220275.236009687, 
    -1887303.21203001,
  
    14941.1540230384, 
    -3206674.8261899,
  
    36843.3319172153, 
    -1957646.01048094,
  
    403506.372278702, 
    -1074722.26073894,
  
    687860.618424752, 
    -2126387.54230178,
  
    447138.947217192, 
    -2286068.61962964,
  
    214315.007728907, 
    -1419951.45431663,
  
    183825.364703231, 
    -1492562.20256775,
  
    256007.951577538, 
    -1795432.27517146,
  
    483331.984120874, 
    -1875917.63550577,
  
    -23288.5861640593, 
    -2502971.01821319,
  
    110328.512350628, 
    -3081727.5389567,
  
    299541.308187916, 
    -2552570.37853665,
  
    -240841.075491053, 
    -1283495.72253156,
  
    -104901.986266784, 
    -3120661.60396672,
  
    198250.896643734, 
    -1672263.88492333,
  
    -531890.354210781, 
    -1346113.57838758,
  
    -187389.154827117, 
    -1666925.33498539,
  
    -38340.4357512889, 
    -1920306.1139364,
  
    570620.098137623, 
    -1465638.38163872,
  
    -96329.9256664722, 
    -3173382.02329799,
  
    -342046.480291845, 
    -1212507.64744466,
  
    243699.712293553, 
    -1936281.7107618,
  
    299010.940748785, 
    -1199752.72756303,
  
    237738.733346825, 
    -2250121.3319434,
  
    428235.649317861, 
    -1127439.93544703,
  
    947.891199243349, 
    -1463679.74414594,
  
    610036.714344292, 
    -2189061.54399711,
  
    6969.6764366514, 
    -2646126.99018783,
  
    402224.292585647, 
    -1422074.07854677,
  
    397357.624628959, 
    -2531551.50203985,
  
    -60593.8512409515, 
    -2638291.90907986,
  
    209338.830872271, 
    -976075.65900022,
  
    280797.439293299, 
    -1907124.24940589,
  
    418216.100988187, 
    -1187981.20956433,
  
    245177.10254334, 
    -2222019.52171563,
  
    193906.505568672, 
    -2548555.10125537,
  
    101715.661428636, 
    -3117391.65731137,
  
    -169798.832739596, 
    -3076899.31983936,
  
    -334216.30692454, 
    -1231997.78185951,
  
    -55993.6452001093, 
    -1664331.30790652,
  
    448831.687150133, 
    -2534559.73959677,
  
    -300544.722643389, 
    -1749214.79726437,
  
    18859.5304889376, 
    -2050266.89541072,
  
    244323.397786818, 
    -920561.608851949,
  
    -346292.343280648, 
    -1450624.62755234,
  
    30452.0013550163, 
    -2490236.00377186,
  
    -246179.130939279, 
    -1336427.89950565,
  
    -400809.408137777, 
    -1431926.38286603,
  
    450556.090214757, 
    -1914917.41130006,
  
    46693.9778661625, 
    -2888167.36957394,
  
    23522.1211957058, 
    -2213347.22412871,
  
    496200.513486765, 
    -2329147.5259004,
  
    330796.914608122, 
    -1421060.67758583,
  
    313618.886180773, 
    -1768661.50330917,
  
    405181.821250712, 
    -2495973.11416183,
  
    -216291.343538387, 
    -2656961.86665481,
  
    66634.1620698333, 
    -2914971.06173432,
  
    78262.8944656525, 
    -1938330.86330547,
  
    39021.987806449, 
    -2160766.09527405,
  
    -126206.615073349, 
    -2281136.43798657,
  
    -530312.424304378, 
    -1179649.85817708,
  
    52334.3748927265, 
    -2979701.57250391,
  
    430128.390833397, 
    -1291450.05068483,
  
    243270.090190978, 
    -2011218.67300784,
  
    -81132.6015837808, 
    -2720132.38691849,
  
    -40497.1303303756, 
    -2159101.1643267,
  
    530410.419988327, 
    -2028969.7672829,
  
    -164165.754745542, 
    -2792244.00668917,
  
    -146475.569938332, 
    -1134154.68928043,
  
    -14602.8352656362, 
    -2824471.99521558,
  
    119765.789579924, 
    -3096912.14936765,
  
    -137806.601278902, 
    -2951851.45468741,
  
    394669.252476605, 
    -1713899.39519463,
  
    357848.16750782, 
    -1949507.55953959,
  
    520284.308554611, 
    -2185301.96309277,
  
    106291.297839044, 
    -1458756.94479718,
  
    102843.629129341, 
    -1815499.88503122,
  
    -143710.987631574, 
    -2841499.32162355,
  
    -170702.014966621, 
    -2098452.27206907,
  
    -41413.5185552962, 
    -2484098.71547813,
  
    130885.723200311, 
    -2285578.33237383,
  
    203969.410525308, 
    -2791361.7565488,
  
    102560.466763917, 
    -2616921.31316138,
  
    503377.344504468, 
    -1530335.09838041,
  
    -160370.344103844, 
    -1603651.16239061,
  
    -107968.313839325, 
    -1895870.80503738,
  
    -66521.6427310127, 
    -2896182.91743722,
  
    215281.25075657, 
    -1118007.75036648,
  
    473266.974816781, 
    -1971198.41021712,
  
    -130682.300319232, 
    -2757896.28389815,
  
    167239.839371525, 
    -2212048.38631058,
  
    160111.89350056, 
    -2486921.15193841,
  
    188146.873872859, 
    -1135613.59918867,
  
    169357.445048634, 
    -1695715.97809448,
  
    153924.549843535, 
    -2000180.88300449,
  
    -16794.529911313, 
    -2608513.07233484,
  
    288963.966325924, 
    -1804214.61497997,
  
    -111067.188744155, 
    -1495253.15451074,
  
    -99729.5913759709, 
    -1860515.61241578,
  
    450399.988825826, 
    -1232724.06729202,
  
    363164.848171189, 
    -2289591.51578254,
  
    -103282.513893634, 
    -2515185.92130268,
  
    345617.849167023, 
    -1393041.73859229,
  
    50536.8442926947, 
    -1535580.99351814,
  
    117350.327167588, 
    -1833694.5715006,
  
    434.113136572047, 
    -944565.44979141,
  
    370114.280438719, 
    -2263756.26628487,
  
    -475816.091097466, 
    -1390966.79384841,
  
    56324.224199883, 
    -3204876.64349565,
  
    -47443.919559943, 
    -2363948.86679936,
  
    -189400.579852173, 
    -1158084.70894666,
  
    -315650.811205598, 
    -1217868.17496619,
  
    367356.134154085, 
    -1677540.0643455,
  
    367196.816298893, 
    -1278543.14624241,
  
    -52171.6693578373, 
    -1677837.83834192,
  
    -56966.0574280309, 
    -2052585.44845869,
  
    269218.61902063, 
    -964945.563181623,
  
    84754.8968189761, 
    -1876645.46817286,
  
    -327103.860844562, 
    -1531527.41806732,
  
    116403.477172322, 
    -1949428.9712825,
  
    -124304.644715938, 
    -2562559.42407557,
  
    467252.478124757, 
    -1133034.31433404,
  
    132250.732637375, 
    -1436770.02842123,
  
    -120816.297446775, 
    -2590185.83643603,
  
    267824.952270923, 
    -1465451.38488114,
  
    55244.4626345688, 
    -2678771.01276153,
  
    63573.5602262657, 
    -947074.142586509,
  
    405434.081985681, 
    -1887920.18029751,
  
    62730.5876050181, 
    -2521024.3979237,
  
    231009.200422959, 
    -2514345.44666727,
  
    -272991.384716172, 
    -1361877.60534385,
  
    97443.4623943168, 
    -1669118.63567736,
  
    -522158.118673098, 
    -1339486.48240848,
  
    592741.9776002, 
    -2255056.08377735,
  
    -113094.059756403, 
    -1946820.45458647,
  
    -112252.581167841, 
    -2447696.71863432,
  
    -365122.151773232, 
    -1298671.40476982,
  
    586267.519165562, 
    -1539313.79343725,
  
    323259.857806676, 
    -1928064.67401814,
  
    -88018.2245216926, 
    -2851536.90230649,
  
    219083.642987019, 
    -1141488.40308797,
  
    157200.191935482, 
    -2236295.45295839,
  
    -324291.837874031, 
    -1405038.3583209,
  
    584889.067607627, 
    -2140013.7879798,
  
    432528.647412669, 
    -2525910.79726203,
  
    -132992.796541625, 
    -2612992.4716687,
  
    291823.058696564, 
    -992486.754322225,
  
    202899.537158059, 
    -1919126.79419743,
  
    383277.177289958, 
    -1106450.38949599,
  
    167118.014817678, 
    -2198826.37045754,
  
    -382728.602055846, 
    -1161698.87911687,
  
    104177.520679418, 
    -2035421.26594311,
  
    67896.8433709741, 
    -2722466.84181956,
  
    -168814.57123191, 
    -2126396.09584845,
  
    -110928.799793879, 
    -2769952.90088379,
  
    -331318.804295056, 
    -1370381.45251584,
  
    114842.539365784, 
    -2515392.25815453,
  
    -208662.617526707, 
    -1260316.42060915,
  
    -155694.072918578, 
    -2820116.02043503,
  
    128213.288873482, 
    -2910333.81329865,
  
    -60419.8469374974, 
    -2198937.08527869,
  
    483134.036420086, 
    -1918375.06125258,
  
    -110394.901443547, 
    -3132426.7814998,
  
    244448.602483942, 
    -1435559.24111293,
  
    232218.235773285, 
    -1786750.3191598,
  
    -12773.4545276293, 
    -2887234.66788414,
  
    364.992330430008, 
    -1950333.40809678,
  
    781022.8927781, 
    -2057865.20127708,
  
    -41641.0889904894, 
    -2136799.24064288,
  
    -24061.9296125753, 
    -2282901.23501293,
  
    337542.594638742, 
    -2520317.97541449,
  
    -290159.380721705, 
    -1645540.49625665,
  
    56832.7882083427, 
    -2963152.632535,
  
    347494.875607903, 
    -1224741.47361941,
  
    331730.430411844, 
    -1995826.26405345,
  
    -183143.209969008, 
    -2718534.45123504,
  
    39701.2709757577, 
    -2179541.83328828,
  
    513853.850993073, 
    -2114135.73784625,
  
    -77544.8892301096, 
    -2802076.4265995,
  
    -107320.728784574, 
    -1054719.46165959,
  
    -551280.38990348, 
    -1184067.43176716,
  
    -58202.2341923386, 
    -2969178.63590816,
  
    595126.306572533, 
    -1567043.30808687,
  
    308010.865173318, 
    -1706905.77302438,
  
    279544.500100243, 
    -1968965.36841705,
  
    21878.4565796481, 
    -1472930.52896503,
  
    24472.7477730172, 
    -1832915.42661567,
  
    30463.177912436, 
    -900620.055077571,
  
    641687.561672487, 
    -2169110.19407721,
  
    756990.15767055, 
    -2057661.31156108,
  
    -141969.637752549, 
    -2458590.70612708,
  
    223178.782150433, 
    -2287172.91682098,
  
    25791.3443839633, 
    -2578979.10753811,
  
    516914.766036657, 
    -1637169.82700882,
  
    481509.604998853, 
    -1380353.3882309,
  
    -199709.017409733, 
    -986163.269591,
  
    -79252.1947800798, 
    -1577470.32764235,
  
    -21307.2994393099, 
    -1871956.87054254,
  
    132647.737986745, 
    -1051299.17304335,
  
    -219402.335394835, 
    -2358752.26314788,
  
    -225426.250496743, 
    -956914.722941295,
  
    83424.6747964064, 
    -2441485.6498615,
  
    -137960.08421351, 
    -1032673.69536206,
  
    209747.730259938, 
    -2703080.27133624,
  
    -576623.490108784, 
    -1390291.97618745,
  
    257472.944447896, 
    -1190954.26935854,
  
    83045.8161114442, 
    -1688750.34169849,
  
    72812.7794362073, 
    -2020336.48416837,
  
    209696.501251925, 
    -1832329.96844842,
  
    -175070.618787317, 
    -1877257.86088269,
  
    709190.06373511, 
    -2170220.96547966,
  
    263553.574075478, 
    -1409860.31269674,
  
    -135377.076183886, 
    -968667.868069451,
  
    133425.609501155, 
    -1508828.69147376,
  
    204011.341567678, 
    -1809780.63700543,
  
    89642.9730559876, 
    -919225.338163622,
  
    -76422.5679320631, 
    -2491819.45959612,
  
    -134628.552353257, 
    -2312293.87748981,
  
    -221550.889077205, 
    -1236466.59175894,
  
    260767.04072566, 
    -1674214.42300496,
  
    435774.237497951, 
    -1333286.19477954,
  
    7744.33670879124, 
    -1903960.32059186,
  
    535764.773678147, 
    -1432680.40481328,
  
    195963.625140491, 
    -1941211.93428096,
  
    286061.8616822, 
    -2258416.85946402,
  
    50186.4572877978, 
    -1453588.60007088,
  
    -40394.836375174, 
    -2625392.12142743,
  
    351824.539838607, 
    -1438340.56719462,
  
    428634.307388645, 
    -2495541.18756919,
  
    -17154.482923809, 
    -2653471.57289613,
  
    156763.16662748, 
    -965615.185810345,
  
    327536.179592429, 
    -1899922.72263415,
  
    158548.753654562, 
    -2473929.41518995,
  
    -122714.458895655, 
    -3063851.85127401,
  
    283.045892841227, 
    -1666087.17377436,
  
    -311478.061532497, 
    -1703026.21773101,
  
    -32331.2646589456, 
    -2059174.27270341,
  
    -355276.468584385, 
    -1498770.53327156,
  
    -21767.6946678424, 
    -2474669.65896921,
  
    -387589.458130379, 
    -1382563.5450368,
  
    96580.4924201732, 
    -3138361.55964041,
  
    402820.003061738, 
    -1919847.63481937,
  
    -3320.40485700073, 
    -2874567.63653194,
  
    73887.3011451854, 
    -2221993.30803281,
  
    -336435.730174061, 
    -1485837.97630222,
  
    530892.479383691, 
    -2223618.70669739,
  
    -204445.382114251, 
    -2380143.84289882,
  
    382605.904673856, 
    -1412361.53768695,
  
    366544.696584274, 
    -2527172.83913237,
  
    114278.733397942, 
    -2931612.89690726,
  
    125001.634764784, 
    -1931129.33653386,
  
    350814.879165391, 
    -1030698.83826042,
  
    87419.8345303814, 
    -2175146.20947401,
  
    544512.221508543, 
    -1550518.01060944,
  
    -321676.942955213, 
    -1081469.02470233,
  
    1747.09804765793, 
    -2971228.64681544,
  
    190193.883551823, 
    -2020454.11814743,
  
    -23167.6334820156, 
    -2721040.37262681,
  
    -88616.169925659, 
    -2146836.76481043,
  
    -169968.474475829, 
    -1181815.82732603,
  
    -67003.7660900606, 
    -2822854.19730282,
  
    -185601.303883927, 
    -2941448.16392183,
  
    -144361.812357698, 
    -2184526.94862541,
  
    446664.285555997, 
    -1718095.57040916,
  
    404830.36927056, 
    -1937832.87258523,
  
    538729.479292925, 
    -2137398.97897203,
  
    -87231.5592452419, 
    -3188008.41115563,
  
    158100.288162786, 
    -1450057.80735319,
  
    150817.587820823, 
    -1804839.13475234,
  
    480494.412040165, 
    -2343782.50897071,
  
    -122304.168242545, 
    -2112832.38626947,
  
    16002.8592961329, 
    -2498663.49249649,
  
    73861.4489080644, 
    -2284593.10021864,
  
    147275.395790736, 
    -2639021.12206547,
  
    495777.842487845, 
    -1470361.28701169,
  
    -538629.610358206, 
    -1372966.89568416,
  
    -209041.233852935, 
    -1619359.66176652,
  
    -159964.923849107, 
    -1910219.16687103,
  
    -19981.9836947078, 
    -2921449.52138295,
  
    264861.360382621, 
    -1158032.89655404,
  
    420190.770632687, 
    -1980433.85509891,
  
    -184080.442577845, 
    -2763567.34762882,
  
    119899.672281782, 
    -2199982.50224958,
  
    497865.393065098, 
    -2196379.38812898,
  
    6959.66367039556, 
    -2811668.62279688,
  
    204259.346159002, 
    -2513077.55267671,
  
    -68165.8878889877, 
    -975284.231583968,
  
    65749.6021532679, 
    -3057173.19391973,
  
    221352.477870016, 
    -1699912.15085407,
  
    201240.832950704, 
    -1988423.17974941,
  
    336637.434759881, 
    -1787305.32757417,
  
    -53898.1335832897, 
    -1850330.96820005,
  
    311948.361254564, 
    -2288706.62806372,
  
    -53995.5934061615, 
    -2539545.38449839,
  
    394856.415513614, 
    -1382950.59697248,
  
    658936.235598381, 
    -2230779.85359421,
  
    1865.95454365216, 
    -1551289.49289409,
  
    65353.7171577388, 
    -1848042.93333448,
  
    50014.222762182, 
    -984590.595978531,
  
    536108.357929154, 
    -2183521.20426147,
  
    2996.5210622136, 
    -2393833.72668216,
  
    -170110.393180363, 
    -1111055.58062914,
  
    -327456.0298889, 
    -1263995.18910224,
  
    432928.048935339, 
    -1679585.94698519,
  
    326050.363191721, 
    -1245697.31815372,
  
    -500545.721714682, 
    -1391887.82367358,
  
    -1465.11135396852, 
    -1681930.02731075,
  
    -8298.99342609953, 
    -2040492.08559011,
  
    226136.44632154, 
    -942026.024064978,
  
    130961.23037847, 
    -1860256.55648842,
  
    -250411.645940582, 
    -1894000.1118045,
  
    68667.3900192572, 
    -1954359.19480158,
  
    -173569.895506866, 
    -2546154.36877898,
  
    479206.280653619, 
    -1208135.38877398,
  
    181489.298725911, 
    -1426678.88434625,
  
    602872.242033096, 
    -1483888.97126231,
  
    217425.199781917, 
    -1481717.8759841,
  
    290672.355709742, 
    -1785866.70005516,
  
    464343.579610888, 
    -2496435.4057141,
  
    452172.822284791, 
    -1880718.65352569,
  
    -297926.616450221, 
    -1808778.14535286,
  
    -481835.374784779, 
    -1170313.96346267,
  
    103872.161493733, 
    -3052347.09434852,
  
    272571.69465804, 
    -2537527.62516161,
  
    -253701.1983023, 
    -1314848.47457126,
  
    157888.204374714, 
    -1671004.54526139,
  
    -168840.049997149, 
    -2082927.27946318,
  
    468628.24313141, 
    -1102898.48098747,
  
    -68241.8854049492, 
    -1930911.84970545,
  
    -168361.027401012, 
    -2430971.16351865,
  
    -351444.039124707, 
    -1247597.80366204,
  
    567059.613278995, 
    -1580031.22866844,
  
    275523.770395591, 
    -1932994.89508233,
  
    267040.02322028, 
    -1176446.99860019,
  
    -194305.427069621, 
    -3046773.97395494,
  
    205523.317815922, 
    -2244590.98073722,
  
    608452.46618617, 
    -2147522.09647263,
  
    37881.3708082356, 
    -2659659.27117021,
  
    435824.127664333, 
    -1411229.75196321,
  
    -89553.4284824026, 
    -2628172.13303023,
  
    243034.165570455, 
    -982779.695843019,
  
    249638.277457194, 
    -1911925.26742573,
  
    403916.425781585, 
    -1154612.57303603,
  
    444533.647655765, 
    -1059978.03279585,
  
    -340993.665349916, 
    -1266670.2871622,
  
    -422576.64451645, 
    -1214064.40762794,
  
    -93359.241270923, 
    -1663165.47978454,
  
    -293325.759261181, 
    -1779711.76543737,
  
    52986.7279865339, 
    -2044328.64297787,
  
    -340302.927143807, 
    -1418527.35797716,
  
    64590.4791812392, 
    -2500412.45497789,
  
    -231172.527047259, 
    -1305983.30810188,
  
    57373.7720796011, 
    -3163387.76544532,
  
    79439.0765868044, 
    -2897071.30239012,
  
    -10054.6645329449, 
    -2207583.16892492,
  
    496394.120093371, 
    -2359927.4870028,
  
    -210512.215183757, 
    -2035309.7256378,
  
    -153258.925569315, 
    -3111061.58134997,
  
    296257.590352666, 
    -1426860.10392706,
  
    281058.625138981, 
    -1775897.03073465,
  
    34871.1143456655, 
    -2903876.50331553,
  
    47103.7326295508, 
    -1943131.88132522,
  
    526028.620167079, 
    -1269870.20416479,
  
    6756.75773351178, 
    -2151179.35484302,
  
    -84965.2865969047, 
    -2281848.98306959,
  
    516232.828496924, 
    -1475048.48243924,
  
    51924.3059161248, 
    -3017646.68528249,
  
    -365294.156826223, 
    -1084631.16352977,
  
    519108.602500929, 
    -1704335.21233839,
  
    397074.985234183, 
    -1264766.61980706,
  
    278654.226227719, 
    -2005061.7089351,
  
    -120985.393007846, 
    -2719508.11601207,
  
    -8417.76887750764, 
    -2167277.43131715,
  
    523737.767104033, 
    -2063293.4748131,
  
    -129030.482437913, 
    -2796232.24597347,
  
    -130813.633321993, 
    -1102380.59970509,
  
    19459.2096186394, 
    -2825523.60712485,
  
    360005.898252726, 
    -1711101.94823895,
  
    326526.701862984, 
    -1957290.68146275,
  
    71751.973583595, 
    -1464556.37113851,
  
    71495.2765868097, 
    -1822466.10166501,
  
    615984.997456893, 
    -2122511.38411864,
  
    -80690.7610716041, 
    -2474135.28044434,
  
    168094.104117941, 
    -2286221.19747573,
  
    72316.0015657196, 
    -2601973.35453106,
  
    508648.86951791, 
    -1571936.9559668,
  
    728328.952426814, 
    -2168529.87943576,
  
    -156828.1597259, 
    -956713.1198974,
  
    -127923.084529155, 
    -1593178.82701829,
  
    -73303.9069941015, 
    -1886305.23211826,
  
    -98339.9350284291, 
    -2878908.61281505,
  
    182227.8451576, 
    -1091324.3194888,
  
    508651.110853488, 
    -1965041.44614422,
  
    -95858.2964954499, 
    -2754197.85643401,
  
    198451.291644425, 
    -2220003.44650766,
  
    129984.022580244, 
    -2469071.04560597,
  
    -118669.897541801, 
    -985644.567044742,
  
    216326.491082839, 
    -1158108.43881487,
  
    48065.8291451456, 
    -3031555.39495136,
  
    134694.088111684, 
    -1692918.52894176,
  
    121479.841241201, 
    -2008243.12401267,
  
    257256.979805318, 
    -1815460.75641897,
  
    -129866.003761923, 
    -1867212.51244838,
  
    680808.728323164, 
    -2162585.72547028,
  
    -199465.834554734, 
    -2952285.16405051,
  
    397245.008777324, 
    -2290180.33380906,
  
    -136840.318280989, 
    -2498600.38507862,
  
    541909.637466809, 
    -1931020.98776375,
  
    312792.14016402, 
    -1399769.16862185,
  
    -179728.030431688, 
    -990231.951606335,
  
    440499.808290568, 
    -1085751.35734166,
  
    83025.8570121264, 
    -1525095.18257678,
  
    152014.73155782, 
    -1824128.99883937,
  
    -578419.158800178, 
    -1374764.42994249,
  
    -130927.286871714, 
    -2480380.21684801,
  
    -482642.815304992, 
    -1361282.76570474,
  
    -247183.71103291, 
    -995249.502965907,
  
    -202260.702405346, 
    -1189437.46344136,
  
    -307780.665416732, 
    -1187116.83220882,
  
    86706.6769624042, 
    -884795.139802802,
  
    323996.500220752, 
    -1676187.21924077,
  
    394627.784390712, 
    -1300440.36669088,
  
    -85976.0415324385, 
    -1675109.71072603,
  
    -89410.7662883386, 
    -2060647.68701164,
  
    297368.903663925, 
    -979921.399259812,
  
    53950.6727232911, 
    -1887571.40864947,
  
    552303.403934332, 
    -2294274.38339214,
  
    502182.257664216, 
    -1244566.69524695,
  
    148227.537729392, 
    -1946142.15534507,
  
    245506.769245565, 
    -936507.901014177,
  
    334384.987562486, 
    -2266712.38724255,
  
    -91595.2312117364, 
    -2573451.47907943,
  
    99425.0233763431, 
    -1443497.45599586,
  
    -88296.6938430872, 
    -2604422.01565105,
  
    301424.787349604, 
    -1454607.05829753,
  
    26284.8853932561, 
    -2668651.23671222,
  
    101627.06119512, 
    -954645.283348892,
  
    374274.920149587, 
    -1892721.1983174,
  
    463649.981418986, 
    -1294002.25652528,
  
    96258.9046547646, 
    -2528061.19427234,
  
    39737.9896441961, 
    -3117536.45726445,
  
    202573.997299398, 
    -2498485.23341103,
  
    -75630.0850515942, 
    -3050804.38270844,
  
    58579.2957421194, 
    -1667906.05042515,
  
    554274.479264207, 
    -2262262.93902501,
  
    -142995.509410036, 
    -1957426.19035543,
  
    733665.75215049, 
    -2080625.6525279,
  
    -75459.8110215002, 
    -2458664.39705057,
  
    -374227.583282233, 
    -1332670.76982107,
  
    355083.915908705, 
    -1924777.85833864,
  
    188116.47619594, 
    -1118914.37623168,
  
    124252.48329162, 
    -2230639.38922375,
  
    -329149.395776062, 
    -1437358.20561667,
  
    562909.91447422, 
    -2174044.92481463,
  
    -161952.373783145, 
    -2602872.69561889,
  
    171740.375321951, 
    -1923927.81221723,
  
    369981.359345411, 
    -1075424.27972005,
  
    135817.681254263, 
    -2189526.32367384,
  
    -357568.916219548, 
    -1128635.76487349,
  
    563119.919428029, 
    -1837918.43889837,
  
    -275791.134935152, 
    -1853787.8975713,
  
    138304.718177028, 
    -2029483.01351019,
  
    32362.2097839145, 
    -2721910.21312205,
  
    -136735.209779, 
    -2134572.36283905,
  
    -146118.247121905, 
    -2775370.0838676,
  
    -193461.376558338, 
    -1229476.96511364,
  
    -119687.479716324, 
    -2821227.66765334,
  
    -93996.6326661742, 
    -2193173.03007479,
  
    209909.275773468, 
    -1441358.66771224,
  
    199657.977186518, 
    -1793985.84632722,
  
    481664.613592731, 
    -2397346.20775611,
  
    -44721.5252230499, 
    -2876075.48339402,
  
    -73906.321776526, 
    -2127212.49801475,
  
    15314.5964929433, 
    -2283581.56028621,
  
    -507754.051460656, 
    -1345658.43976443,
  
    -434443.345825394, 
    -1147550.90765773,
  
    -257712.120888973, 
    -1635068.16333941,
  
    -211961.531403833, 
    -1924567.52844656,
  
    26106.8798349735, 
    -2946471.38704067,
  
    314441.470008767, 
    -1198058.04274165,
  
    367114.566448579, 
    -1989669.29998065,
  
    71780.6324285856, 
    -2187718.10027862,
  
    507414.599549899, 
    -2147258.85572099,
  
    -43385.3055505824, 
    -2805953.91415178,
  
    247332.424650828, 
    -2538597.41054637,
  
    -91658.7924263222, 
    -1022945.36962931,
  
    -502188.092304251, 
    -1211689.16495556,
  
    273347.51094943, 
    -1704108.32606867,
  
    248223.034713442, 
    -1976748.49279519,
  
    385552.041380016, 
    -1769955.819461,
  
    -416519.636950531, 
    -1414619.84654078,
  
    -11357.9560433164, 
    -1478511.1848667,
  
    -6875.60476950814, 
    -1839881.64324944,
  
    63769.4057664488, 
    -903025.564449231,
  
    -184472.686533973, 
    -2447808.98164639,
  
    258803.323672307, 
    -2287788.4168838,
  
    -5804.19596503216, 
    -2563363.39715688,
  
    444094.979147161, 
    -1372859.45315571,
  
    -46804.9349473693, 
    -1566997.99472506,
  
    13357.107147899, 
    -1862391.29516833,
  
    -177885.666741753, 
    -2835722.85384302,
  
    99594.329932865, 
    -1024615.74242381,
  
    -150820.209221647, 
    -1064026.45011469,
  
    -339261.248572201, 
    -1310122.20323829,
  
    500215.136310703, 
    -1681685.34112915,
  
    284903.912281592, 
    -1212851.48735198,
  
    49241.4441948753, 
    -1686022.21653761,
  
    40368.0708338896, 
    -2028398.72517649,
  
    177989.514731324, 
    -1843576.10988738,
  
    -205207.031173252, 
    -1883954.76091525,
  
    64219.0919485294, 
    -3220893.89460967,
  
    20931.3026081616, 
    -1959289.4158656,
  
    694806.379598544, 
    -2140661.54268553,
  
    -103867.686585701, 
    -2968626.21787947,
  
    -205859.390526923, 
    -2500833.16070504,
  
    479453.004736546, 
    -1268727.95385011,
  
    230727.862359422, 
    -1416587.74052934,
  
    167025.447034871, 
    -1497984.36463206,
  
    238675.748154906, 
    -1800215.06163111,
  
    48654.86505735, 
    -923876.486333787,
  
    498911.562583887, 
    -1873517.12675384,
  
    -40999.9143244081, 
    -2499253.83127519,
  
    -234411.014085432, 
    -1267819.34651171,
  
    218905.860181269, 
    -1672908.32997283,
  
    463205.205331772, 
    -1355183.41277297,
  
    -23059.8873868777, 
    -1914886.2610684,
  
    559001.656651133, 
    -1454652.38936358,
  
    -114070.99288051, 
    -3173029.48033478,
  
    683692.724382405, 
    -2086407.20307745,
  
    227787.683242532, 
    -1937925.11860152,
  
    253846.44369631, 
    -2252886.50851595,
  
    17360.7455717318, 
    -1460316.02790358,
  
    610828.837324828, 
    -2209831.26911574,
  
    -8486.16816511727, 
    -2639360.85066607,
  
    385424.374917288, 
    -1427496.24061104,
  
    407783.184816516, 
    -2519548.06478736,
  
    -46114.0601652121, 
    -2643351.79684661,
  
    191971.19320824, 
    -972620.186403987,
  
    296377.017756326, 
    -1904723.740654,
  
    425462.079047622, 
    -1204889.8754059,
  
    -567947.587237755, 
    -1151585.98768174,
  
    85715.6650892307, 
    -3124063.46338222,
  
    -154104.039821612, 
    -3072550.16347891,
  
    -37310.844709677, 
    -1664914.22170948,
  
    355428.872742031, 
    -1493850.29804064,
  
    337521.080247462, 
    -1538871.42670864,
  
    413733.857393838, 
    -2204422.52172948,
  
    294756.534747456, 
    -2020260.65439668,
  
    366420.47447029, 
    -1532430.35009665,
  
    134407.484494347, 
    -1913182.47184143,
  
    -87245.9894877849, 
    -2099131.63766289,
  
    -94221.429748457, 
    -1630390.59182323,
  
    19531.1671325101, 
    -2067884.53552615,
  
    -34222.5439729805, 
    -2930599.27934322,
  
    126410.541230812, 
    -1681737.79715941,
  
    -250526.417734201, 
    -1550146.02852206,
  
    497722.004267635, 
    -2118213.12068377,
  
    -51923.5305934056, 
    -2672305.91335474,
  
    129478.546879627, 
    -1609437.2240735,
  
    510684.731476275, 
    -1998544.84834565,
  
    -183309.716442127, 
    -3018703.58915793,
  
    70571.8553429148, 
    -2303291.9004038,
  
    -213801.867443067, 
    -1044449.11013836,
  
    16379.7588393515, 
    -2003399.74014378,
  
    125604.037983466, 
    -1295859.86855395,
  
    -7470.25666767299, 
    -2673159.19876895,
  
    363265.075498708, 
    -1341266.74869248,
  
    236776.641340142, 
    -2370324.55621741,
  
    292113.962360538, 
    -2134276.09315862,
  
    13516.675647145, 
    -2628293.49117986,
  
    151986.020441632, 
    -2554346.58621297,
  
    -27550.810843926, 
    -1778820.55483791,
  
    103629.440890898, 
    -2162138.78828238,
  
    128598.144142173, 
    -2266631.76273907,
  
    159713.015244405, 
    -1024817.45528562,
  
    -317823.867936638, 
    -1617752.02912948,
  
    449677.164625601, 
    -1992053.30760512,
  
    -128508.511598591, 
    -2094910.70677904,
  
    367619.139796618, 
    -1116427.76642336,
  
    526291.665272025, 
    -2125767.35963667,
  
    60065.7270186022, 
    -1105320.02332194,
  
    -116010.380070206, 
    -2367680.43311392,
  
    124911.011373848, 
    -2502926.87509618,
  
    -120100.183976883, 
    -1627302.66437483,
  
    17477.2177648095, 
    -1717076.79386368,
  
    275463.113523234, 
    -1262944.62281326,
  
    -15006.8450097206, 
    -2576793.07784176,
  
    324604.03040553, 
    -2068180.29275127,
  
    -79895.7600063566, 
    -1741349.1115891,
  
    125793.590831948, 
    -2133800.29822904,
  
    -137325.122250525, 
    -2628693.99498834,
  
    -135620.133020713, 
    -1323429.18601639,
  
    148497.903481922, 
    -2430375.36019392,
  
    104847.464060327, 
    -1902746.03160242,
  
    -349946.82254437, 
    -1090552.95086296,
  
    164086.258515934, 
    -1864373.42052164,
  
    -14521.5166294834, 
    -2772100.62137136,
  
    127313.106137732, 
    -2304148.24309085,
  
    244554.878856359, 
    -2153239.19874023,
  
    129767.806110318, 
    -892892.236150582,
  
    -86471.0706210469, 
    -2383352.1015983,
  
    -294619.76349246, 
    -1101938.98819075,
  
    53713.5449677728, 
    -1061509.37953705,
  
    -169550.698789784, 
    -2162670.0061488,
  
    -279141.365553332, 
    -1213053.46557425,
  
    192695.591508399, 
    -1179493.80033522,
  
    -24797.1199010796, 
    -2262229.08860702,
  
    -214171.606637169, 
    -1862834.6067314,
  
    -275859.5242751, 
    -1489413.25503952,
  
    155219.244839712, 
    -1612629.06872128,
  
    -85130.1970991362, 
    -1792244.95920811,
  
    184512.04699976, 
    -2450229.66318779,
  
    527664.530562995, 
    -1446468.98300822,
  
    -129519.690109271, 
    -2123702.3759108,
  
    -44793.6217871247, 
    -1055928.61444978,
  
    449176.849371941, 
    -1437751.62662047,
  
    -26714.7159117395, 
    -1595317.7094975,
  
    105675.969362104, 
    -1965194.6139386,
  
    166090.017188163, 
    -2075648.52385743,
  
    -344482.854902563, 
    -1167186.67404851,
  
    41771.8849762063, 
    -2855104.67676035,
  
    230655.942358725, 
    -1249522.66435481,
  
    484020.060558395, 
    -1986227.93931313,
  
    83740.0870438672, 
    -1860270.37139919,
  
    -163209.204862947, 
    -2974121.80107097,
  
    76942.8635697521, 
    -1334118.7854879,
  
    414888.407571542, 
    -1794357.31835584,
  
    118028.849710367, 
    -1761023.31598104,
  
    -101417.478400956, 
    -1760394.09886321,
  
    135885.696811887, 
    -1985183.88799928,
  
    -74663.3317180911, 
    -2247050.07235575,
  
    -183835.763421706, 
    -2140986.19212607,
  
    438585.923644013, 
    -1360228.98590885,
  
    655986.354697357, 
    -2115195.22788843,
  
    7618.59673554091, 
    -1588483.25400596,
  
    160026.707700746, 
    -1254038.10309214,
  
    -63855.2005084678, 
    -1385612.1513932,
  
    -69973.1259149521, 
    -1050095.53246778,
  
    207292.719902569, 
    -1010213.22855497,
  
    344159.584874136, 
    -1726873.68506959,
  
    190952.902120091, 
    -1261345.14194011,
  
    7089.15550003367, 
    -1446494.28501419,
  
    120366.000436317, 
    -2118094.32402795,
  
    -203976.772176464, 
    -1430412.83376936,
  
    -5846.88016432955, 
    -3063800.14274786,
  
    71539.9761583662, 
    -1061262.59924972,
  
    301200.01194825, 
    -1386856.55639395,
  
    -144186.3777954, 
    -1383947.8084962,
  
    44648.5508720358, 
    -1104082.13095393,
  
    443382.212766692, 
    -2385299.24772519,
  
    120279.472301642, 
    -2248172.3767743,
  
    -118932.390456188, 
    -1704971.27769198,
  
    -127764.625612486, 
    -1529755.2648849,
  
    54883.8051878682, 
    -1720616.96659444,
  
    119700.859195245, 
    -2840931.23283704,
  
    214922.377887079, 
    -1356926.3442839,
  
    -167445.373393934, 
    -1994985.79962821,
  
    -88378.2668647419, 
    -2540369.83250689,
  
    -61650.5917848601, 
    -2094677.95024414,
  
    -104144.468402464, 
    -2610731.85112339,
  
    -90409.6581521533, 
    -2162282.18828797,
  
    293320.516733886, 
    -1948212.6466708,
  
    383904.86566444, 
    -1205815.88642772,
  
    -91362.8524150625, 
    -1261815.38928677,
  
    -142671.211465232, 
    -2595909.89015803,
  
    -44174.3633982392, 
    -1361439.36425782,
  
    539091.68749263, 
    -2084978.34192903,
  
    328610.348518972, 
    -1746079.51450525,
  
    244903.355833003, 
    -1895174.29376504,
  
    -36691.5446639741, 
    -1011478.26313701,
  
    -17198.4451586121, 
    -1696770.41573654,
  
    -151078.983048065, 
    -1347043.69572709,
  
    363727.385125713, 
    -1813311.14283387,
  
    464234.247627182, 
    -2345328.93062174,
  
    387013.137598283, 
    -2414293.18244738,
  
    23597.5468826233, 
    -1931675.03539072,
  
    -74275.0458758787, 
    -1986341.56599481,
  
    445726.13129692, 
    -1661391.4707731,
  
    501940.548450434, 
    -1930619.73151649,
  
    41711.7407388636, 
    -3192347.31487828,
  
    -354745.506543279, 
    -1196647.56521125,
  
    51365.9674373683, 
    -1630127.64819558,
  
    -14068.1135948399, 
    -2424034.0661133,
  
    297404.646032374, 
    -1612996.89661496,
  
    13926.9867443121, 
    -2958850.01964114,
  
    451525.227137983, 
    -1817032.22624988,
  
    38146.7668012784, 
    -2128718.99450631,
  
    -125937.49032026, 
    -1236170.38458798,
  
    411209.312571803, 
    -1853568.84285074,
  
    507478.158249951, 
    -1780770.24332781,
  
    230045.082822838, 
    -1769382.68663555,
  
    67894.6831057842, 
    -2059333.16396757,
  
    -172981.958258116, 
    -1865980.03557641,
  
    90567.4646658443, 
    -1736905.44847744,
  
    223568.283670922, 
    -1203406.62837193,
  
    -101983.308989316, 
    -1443721.24659755,
  
    -30014.1391221715, 
    -1859033.51077198,
  
    2961.13509942596, 
    -1850825.38827543,
  
    -187988.124798518, 
    -1576589.92745652,
  
    183737.26562071, 
    -1975828.27615092,
  
    -169286.045460385, 
    -1000842.39019381,
  
    36480.7319925061, 
    -3051554.51603057,
  
    253008.844171253, 
    -1734878.78450824,
  
    -93936.9886551359, 
    -3088631.43299373,
  
    -57910.3339590008, 
    -1333140.89685653,
  
    -203072.41837745, 
    -2900571.29059809,
  
    -21989.783818482, 
    -2838139.28380015,
  
    62521.8018337669, 
    -2576888.05069331,
  
    -13055.1061670799, 
    -1516295.50495514,
  
    35537.5622669968, 
    -1843164.55867631,
  
    460402.911292416, 
    -1956936.33697549,
  
    119845.619365881, 
    -1708426.84844271,
  
    424749.637012507, 
    -2230768.89054916,
  
    63367.036070679, 
    -2931031.58796166,
  
    -174800.94747543, 
    -2256247.76134976,
  
    -155604.699787755, 
    -1733941.98504194,
  
    143843.578250353, 
    -2250412.63072641,
  
    -158203.580344285, 
    -2589803.44387565,
  
    255956.126665011, 
    -1051304.97761302,
  
    -32899.7597347711, 
    -2532721.43370964,
  
    240564.278294323, 
    -1319313.6525612,
  
    285116.249593761, 
    -1008004.94225944,
  
    71204.2286771756, 
    -1433569.9765641,
  
    89403.7566771581, 
    -1632756.44969333,
  
    -255631.82171351, 
    -1273481.57329539,
  
    -26873.0347829899, 
    -2125108.9459922,
  
    -67960.7426959069, 
    -3140704.91688041,
  
    437997.396477938, 
    -1729759.23080674,
  
    -14817.6565252354, 
    -2319532.21179859,
  
    -154426.808855966, 
    -1479557.54469947,
  
    318943.734629572, 
    -2491723.42936294,
  
    193209.405793779, 
    -1609461.06825449,
  
    162688.398345275, 
    -2457191.90840438,
  
    -263767.166557591, 
    -1476877.85904245,
  
    479890.822306443, 
    -1462161.28057055,
  
    32965.9919189313, 
    -2528958.22271347,
  
    46417.2471871207, 
    -2250393.98755674,
  
    324915.196949415, 
    -2229025.18616339,
  
    -328621.277292241, 
    -1555637.54426638,
  
    391372.581196468, 
    -2353849.39469517,
  
    305057.144777403, 
    -2528922.8015156,
  
    378257.106877861, 
    -1133939.93948177,
  
    74796.2328029594, 
    -973981.16690414,
  
    264963.725131714, 
    -1234931.32134835,
  
    446815.015481348, 
    -2256773.56392962,
  
    343217.340526221, 
    -1656469.33360646,
  
    353577.653178569, 
    -2229075.80742155,
  
    -288647.785768511, 
    -1738875.2067517,
  
    415954.995109589, 
    -1231737.22604707,
  
    379120.016379473, 
    -1733105.22708532,
  
    -300351.100049786, 
    -1118634.37980141,
  
    203527.781808774, 
    -962271.5378964,
  
    481637.494558538, 
    -1640857.64630264,
  
    47660.4429491012, 
    -2924543.05840613,
  
    297286.751412914, 
    -2334775.31500524,
  
    -44705.3847209393, 
    -3089768.04278716,
  
    474498.272547054, 
    -1442393.72668822,
  
    205623.725994959, 
    -2156286.3992483,
  
    316833.5744338, 
    -1277857.1754933,
  
    231305.326165569, 
    -1015065.09893418,
  
    293906.408601469, 
    -1918037.61394831,
  
    200043.575536941, 
    -2174093.31363477,
  
    -229715.512817201, 
    -1084999.47090455,
  
    -232355.634168386, 
    -1551503.73898993,
  
    122699.690268685, 
    -1343868.79283148,
  
    350397.929451094, 
    -1554921.49549749,
  
    318834.781803247, 
    -1542050.04668407,
  
    194006.215191451, 
    -2473843.92705237,
  
    311214.910776281, 
    -2105288.04411159,
  
    -363888.439906159, 
    -1226438.2530133,
  
    276903.010677481, 
    -2180871.95412809,
  
    343309.034537653, 
    -1300638.19413683,
  
    344911.816549771, 
    -1056369.04595074,
  
    -56715.0142323877, 
    -2381798.59250253,
  
    -185645.415394105, 
    -2222422.55978497,
  
    -146746.767483356, 
    -2863157.98537946,
  
    -106445.039387289, 
    -2262018.75276428,
  
    285884.161211394, 
    -1123310.1044455,
  
    -18155.0003871154, 
    -3086176.51379041,
  
    -22858.1799812265, 
    -2953650.06935816,
  
    454180.852999204, 
    -2066169.78261844,
  
    -275598.460846253, 
    -1270768.36754373,
  
    198344.486882346, 
    -1823567.62504375,
  
    459925.083276316, 
    -2277379.01253003,
  
    -114862.589293503, 
    -2684691.76173705,
  
    303465.550686855, 
    -1266587.18222826,
  
    253301.216321092, 
    -1331697.63733223,
  
    186137.241694357, 
    -1713862.85518005,
  
    339452.14983023, 
    -1880456.17199247,
  
    -66262.8331878217, 
    -1708677.61846454,
  
    -224175.555052987, 
    -3001081.7051218,
  
    -160278.145769936, 
    -2617055.78818607,
  
    -151839.779044989, 
    -1321118.49240913,
  
    -54493.3195120531, 
    -2016250.41233524,
  
    119245.283299903, 
    -2049093.3413829,
  
    456152.802403792, 
    -1384928.61617873,
  
    -438.427166978821, 
    -2071866.01558386,
  
    88698.1202684728, 
    -2424162.61780059,
  
    -278372.307862452, 
    -1572713.07765588,
  
    -174387.357032034, 
    -2740936.68390878,
  
    116483.021063168, 
    -2763686.94808897,
  
    409760.921481733, 
    -1951507.41038638,
  
    89343.1457191578, 
    -2846084.86798008,
  
    -122294.067556676, 
    -2886185.01436422,
  
    -134380.764582705, 
    -2334283.67266635,
  
    189940.674225242, 
    -1198064.9055637,
  
    -211283.730906701, 
    -1692364.92749325,
  
    -91035.4499422129, 
    -2921331.77066982,
  
    117787.075116522, 
    -2662513.28748103,
  
    292243.789679542, 
    -1257629.22967683,
  
    -81880.8169555212, 
    -1524371.35982776,
  
    205299.841887277, 
    -2338836.33851254,
  
    -73367.8889018789, 
    -2074265.55150041,
  
    137742.808277822, 
    -2065642.4643879,
  
    506375.410068381, 
    -2084215.60141067,
  
    -109698.360281239, 
    -1341272.96395373,
  
    -152917.383380104, 
    -3058704.71085897,
  
    175912.498973849, 
    -2758138.1090344,
  
    176181.189668238, 
    -2128769.67222463,
  
    282261.374857045, 
    -1147552.79955661,
  
    -232299.509530769, 
    -1380110.79311973,
  
    87599.4367742583, 
    -2467320.99375597,
  
    251612.380147915, 
    -2134824.83101332,
  
    381680.403672211, 
    -1369139.5226434,
  
    -395699.889495199, 
    -1258847.34891394,
  
    13653.6763361238, 
    -3010703.84547451,
  
    296362.584331991, 
    -1691244.35712852,
  
    379001.278339515, 
    -1965535.85287745,
  
    268992.636448179, 
    -1483078.26432645,
  
    125445.090546856, 
    -1407553.7515092,
  
    14866.7590667106, 
    -2918229.99781786,
  
    77142.3517676103, 
    -2121532.94621603,
  
    -244223.141534039, 
    -1614194.01335586,
  
    -122843.38184465, 
    -3094499.14221781,
  
    390847.092910007, 
    -2484364.15465036,
  
    -313930.514155868, 
    -1430970.65887645,
  
    -268280.278785989, 
    -1227528.75328551,
  
    -89476.7072020586, 
    -1330460.1830812,
  
    -71251.3269302032, 
    -2981869.05453501,
  
    -76662.8289172998, 
    -2702321.7442166,
  
    -363930.230554104, 
    -1488275.25213828,
  
    -275255.31972269, 
    -1187197.58778918,
  
    -108741.96784103, 
    -2174443.54755219,
  
    -291237.534614695, 
    -1843793.96803146,
  
    231320.802853639, 
    -2650975.38582388,
  
    223001.405045426, 
    -1262230.06934698,
  
    -79181.019509342, 
    -1111971.11699136,
  
    494825.985653573, 
    -1587033.3820294,
  
    76936.4769338188, 
    -2617830.08821933,
  
    -23944.2570950155, 
    -1130391.8429958,
  
    2012.85994273114, 
    -1734273.52686279,
  
    108716.190564755, 
    -2302609.44809325,
  
    -104644.129247395, 
    -1814403.20821019,
  
    288768.18736912, 
    -1873693.27382596,
  
    287748.723365184, 
    -1985087.81194188,
  
    103702.328505502, 
    -2493634.87581754,
  
    -205000.918886239, 
    -1153457.20256315,
  
    360920.368159038, 
    -2331933.24265301,
  
    -301994.929763175, 
    -1673048.0226729,
  
    117894.863967295, 
    -1379403.14617331,
  
    -154534.029574074, 
    -1255271.55748853,
  
    -89577.9119630203, 
    -1076933.23025609,
  
    246942.117712631, 
    -1882182.81694782,
  
    -20030.5567002284, 
    -2685789.54825575,
  
    164439.827877841, 
    -1349143.81122584,
  
    -136713.088701457, 
    -1252989.85549298,
  
    -210490.674328605, 
    -1473561.69206263,
  
    86778.8517092792, 
    -1984104.93647229,
  
    -49793.3166826897, 
    -1004709.26894805,
  
    -3666.94960198311, 
    -1746209.5080017,
  
    -145483.472043142, 
    -1369616.79891298,
  
    218665.321247851, 
    -2373567.82880091,
  
    432909.751494444, 
    -1470413.99437618,
  
    -132813.046471422, 
    -2037670.0524306,
  
    -100568.815506238, 
    -2031258.05640831,
  
    53249.2968307528, 
    -1810474.58737932,
  
    -42586.6800525433, 
    -2187579.79923706,
  
    211260.630873009, 
    -1595217.06750612,
  
    -183194.132672527, 
    -2066199.58013294,
  
    -194775.473669214, 
    -1032688.19955559,
  
    47353.353044967, 
    -2761109.12380657,
  
    294641.171544864, 
    -1515020.6963856,
  
    18982.8633001478, 
    -2338877.43631368,
  
    449579.804123108, 
    -1761649.19396286,
  
    39178.7089873201, 
    -1439999.96285468,
  
    256216.680126132, 
    -1505401.58222843,
  
    -125280.791758443, 
    -2171159.48359697,
  
    201112.25065489, 
    -1762161.70844269,
  
    79075.7036974311, 
    -2937509.98082226,
  
    -155277.813131346, 
    -1567748.15427675,
  
    -381402.829893873, 
    -1297726.13312648,
  
    171482.699726502, 
    -1396050.82886475,
  
    -219281.884357805, 
    -1318208.40229578,
  
    -45478.5944812882, 
    -1517254.30426351,
  
    -65499.0920304169, 
    -1628832.43834525,
  
    -345741.324007934, 
    -1143507.80178576,
  
    407249.603987475, 
    -2345857.32819719,
  
    -123854.051711402, 
    -2903533.59473213,
  
    -263528.844357239, 
    -1602438.08704104,
  
    467837.874770855, 
    -2265894.22695076,
  
    -267098.497292442, 
    -1309116.08122412,
  
    107926.456441782, 
    -1852340.06370907,
  
    -249129.335710136, 
    -1462148.32098647,
  
    395420.555158073, 
    -1856877.7562305,
  
    34737.0891577707, 
    -1797437.65816097,
  
    -48528.540149854, 
    -2774290.40221756,
  
    -153011.875130401, 
    -2165954.06764903,
  
    455821.652898184, 
    -2244144.94856146,
  
    164585.722935459, 
    -1783404.02075694,
  
    -9910.59556141154, 
    -2343688.53892419,
  
    168665.937946549, 
    -2632186.10297812,
  
    -172356.503845984, 
    -1780539.42218621,
  
    648170.339032156, 
    -2103068.45297712,
  
    -121952.407455507, 
    -2633146.16143967,
  
    357755.011596115, 
    -2381850.11858776,
  
    34302.1851412301, 
    -2432415.52953142,
  
    -54523.8417470418, 
    -2937564.58113644,
  
    84907.5426400233, 
    -1348759.49028986,
  
    63849.0705024061, 
    -1514596.08881852,
  
    78770.4232440609, 
    -1478335.53354652,
  
    8077.12221163948, 
    -1935096.36440088,
  
    171522.620721408, 
    -1632079.05413549,
  
    397176.222717225, 
    -1453559.28948153,
  
    -427906.224287833, 
    -1337340.80754741,
  
    -322789.354512506, 
    -1462806.95854411,
  
    253160.983950889, 
    -2373708.58704464,
  
    39474.0864923108, 
    -2010453.65304401,
  
    -205300.577264166, 
    -1938894.65891163,
  
    10873.8590142338, 
    -2245742.69085485,
  
    481775.465932306, 
    -1480928.80541057,
  
    411320.127531687, 
    -2245153.56598721,
  
    646500.506473352, 
    -2200257.35962717,
  
    346406.280570829, 
    -1199381.8331242,
  
    -82976.1284327633, 
    -2320462.73360702,
  
    -28220.5298926591, 
    -2028531.42422447,
  
    473427.019242136, 
    -1527209.36040634,
  
    246939.879144196, 
    -1571107.5892757,
  
    203860.36289865, 
    -1869983.24542802,
  
    -9630.31431637313, 
    -1591902.13362554,
  
    242059.395351714, 
    -1272738.98078246,
  
    467484.487475805, 
    -1986288.41909544,
  
    136234.642526118, 
    -1198370.20074003,
  
    -73933.4946347157, 
    -2372683.48950884,
  
    352580.385168481, 
    -1865232.54901381,
  
    -30966.3493838174, 
    -2223022.80351119,
  
    -262631.154671676, 
    -1727872.72757938,
  
    304441.760120302, 
    -1870257.7248063,
  
    -266330.591164424, 
    -1132334.4391012,
  
    552076.586464475, 
    -2224430.42082374,
  
    229554.609615567, 
    -2440570.71530277,
  
    175250.337725087, 
    -1478394.07263828,
  
    46678.4577181124, 
    -2570249.4446233,
  
    305342.837181208, 
    -1723249.14658831,
  
    347525.732518282, 
    -2485800.04616317,
  
    248658.233256186, 
    -2591269.89965353,
  
    331141.909440281, 
    -2013104.92551801,
  
    232252.469193331, 
    -2085036.79863851,
  
    286440.118936282, 
    -1372147.01970567,
  
    -91169.0779823501, 
    -1923226.11103488,
  
    135733.651519868, 
    -1595919.04522041,
  
    191704.753053346, 
    -2137074.09820603,
  
    21904.072979234, 
    -2383560.09133585,
  
    165698.275079008, 
    -949388.562795662,
  
    43671.5156735902, 
    -3007684.5919949,
  
    354210.067552038, 
    -1475079.68211497,
  
    333544.7166051, 
    -1520389.90962225,
  
    428816.803099193, 
    -2197624.1626506,
  
    -41258.0249867365, 
    -1950677.40404341,
  
    363410.99008109, 
    -1513030.3008896,
  
    117951.473100163, 
    -1882291.75702926,
  
    -93915.8245709322, 
    -2085091.20761592,
  
    279769.413556385, 
    -957997.589900603,
  
    -93790.3366081864, 
    -1646778.03716042,
  
    101930.801479024, 
    -1537521.08665429,
  
    -245474.106347009, 
    -1565035.98939311,
  
    378981.538513851, 
    -2002998.67193955,
  
    -48965.7894246319, 
    -2657564.67163529,
  
    500821.887220223, 
    -1983332.38887694,
  
    -167660.555673871, 
    -3008838.92618034,
  
    67282.2615197344, 
    -2321990.69813386,
  
    -201271.484753514, 
    -1057181.6338851,
  
    20262.7359092831, 
    -2017914.79371946,
  
    130380.35830186, 
    -1278926.35052672,
  
    -4066.01018118972, 
    -2704686.78561301,
  
    369147.482639242, 
    -1324008.41889789,
  
    241181.977418781, 
    -2353817.32938443,
  
    294771.959170351, 
    -2117864.3904868,
  
    -328886.522866785, 
    -1332948.27052966,
  
    -28801.068908471, 
    -1762684.50572024,
  
    102052.108139939, 
    -2053142.85715428,
  
    333354.033225063, 
    -1913171.99440628,
  
    -446004.39651152, 
    -1140588.95775218,
  
    154520.842746551, 
    -1044437.76209494,
  
    -288365.84058639, 
    -1631192.69712837,
  
    511472.776014366, 
    -2051016.6041588,
  
    351461.50104866, 
    -1126723.48891869,
  
    501099.072775769, 
    -2101529.44568887,
  
    -107674.964787645, 
    -2350441.13786531,
  
    134979.48532088, 
    -2490461.48686971,
  
    -116058.398299098, 
    -1644933.10759825,
  
    -128421.121514193, 
    -1610132.2467734,
  
    16457.1450215581, 
    -1700185.44262022,
  
    272316.180603775, 
    -1279642.33463369,
  
    322859.059024698, 
    -2085896.92603034,
  
    -78375.6892046018, 
    -1757908.95989902,
  
    123757.417145083, 
    -2150777.84943404,
  
    -141858.065269542, 
    -2645122.60580293,
  
    -124696.935808789, 
    -1336485.02869474,
  
    146100.377451539, 
    -2448012.11512715,
  
    102502.978052041, 
    -1886969.26591577,
  
    -331500.356086804, 
    -1118439.51432003,
  
    166036.499243379, 
    -1879547.66004934,
  
    -9298.02711426233, 
    -2791258.37328156,
  
    123740.48881712, 
    -2322718.15135277,
  
    244710.435520886, 
    -2170434.28064718,
  
    -97529.7451902157, 
    -2398063.0629149,
  
    -265570.437597887, 
    -1101722.84167833,
  
    36042.6406558039, 
    -1064007.97849701,
  
    -5016.89125887652, 
    -961665.276291736,
  
    -208140.070754362, 
    -1232942.1727137,
  
    197499.199005855, 
    -1163203.80485653,
  
    -226187.99704538, 
    -1853948.75274183,
  
    -268245.28239184, 
    -1504889.68090973,
  
    154351.242381071, 
    -1593644.12339296,
  
    -85247.3993188051, 
    -1776014.40677904,
  
    178953.349504894, 
    -2466219.81692179,
  
    30252.4692170887, 
    -2703421.39488132,
  
    434100.527357948, 
    -1427201.77180952,
  
    -24744.720481814, 
    -1612414.1465219,
  
    110860.49034487, 
    -1979316.84629994,
  
    168227.282613936, 
    -2058276.55061312,
  
    -356951.581766272, 
    -1156407.04880415,
  
    35897.201053335, 
    -2869369.40181186,
  
    233931.320884416, 
    -1232143.41253268,
  
    494773.146299992, 
    -2001257.4684091,
  
    -150356.022385614, 
    -2962853.47501436,
  
    80765.2077677089, 
    -1317051.66659014,
  
    408378.036623854, 
    -1779277.43909978,
  
    118191.835672779, 
    -1778021.13532115,
  
    -101709.627107885, 
    -1743064.40984404,
  
    121667.080318959, 
    -1962967.63705069,
  
    -79726.2424623726, 
    -2264152.04969468,
  
    -169758.295167242, 
    -2112424.18789935,
  
    10556.5785333121, 
    -1607478.78963975,
  
    164043.87387233, 
    -1237120.31615562,
  
    -53054.6872697138, 
    -1398623.41706702,
  
    216887.135791162, 
    -994580.074800396,
  
    345644.952548055, 
    -1744044.14744601,
  
    195181.832558402, 
    -1244139.02651826,
  
    -186815.043054887, 
    -1185731.98051039,
  
    -215418.566128849, 
    -1417704.7658432,
  
    4468.65609330514, 
    -3078743.85818848,
  
    306020.740559985, 
    -1370580.22766571,
  
    -132831.68518462, 
    -1397260.20756937,
  
    463453.104183242, 
    -2377208.18186612,
  
    58693.8779426751, 
    -2397902.70044657,
  
    -119356.401952598, 
    -1688676.43162858,
  
    -127804.239727899, 
    -1545611.15535376,
  
    52062.6234638594, 
    -1703319.59169506,
  
    117764.448558081, 
    -2857176.66916236,
  
    210667.321076157, 
    -1373523.55030342,
  
    -131801.923110382, 
    -1851087.81594333,
  
    -90000.5973803412, 
    -2557053.05625299,
  
    -67778.4569097129, 
    -2110945.22290195,
  
    183424.00167304, 
    -1152002.98063096,
  
    -9417.57223620058, 
    -1449785.86756765,
  
    316549.799964531, 
    -1753572.25225348,
  
    401314.450897221, 
    -1196766.53995381,
  
    -101473.517365892, 
    -1248117.3013809,
  
    -55309.7862715539, 
    -1347794.65850119,
  
    338528.083227316, 
    -1407158.98582718,
  
    358334.843690165, 
    -1797416.65183203,
  
    503871.87970955, 
    -1651775.06791053,
  
    -476485.788779179, 
    -1243353.80323168,
  
    516762.544977856, 
    -1945450.82207978,
  
    235661.236828563, 
    -1653711.20065129,
  
    47844.6579077996, 
    -1611685.47348197,
  
    -5535.79613730236, 
    -2408933.89762528,
  
    295726.948746057, 
    -1592915.68119259,
  
    -200122.845240878, 
    -1901176.48776782,
  
    447319.209773288, 
    -1801147.16916215,
  
    37709.1599812302, 
    -2112695.44373532,
  
    -114929.742019853, 
    -1249759.02180417,
  
    416122.632570827, 
    -1869580.57851615,
  
    227871.932327411, 
    -1752015.05385323,
  
    65739.0430297559, 
    -2077306.80955909,
  
    88060.2493853987, 
    -1720853.74695015,
  
    226805.128915063, 
    -1186231.83999753,
  
    -89556.7167371838, 
    -1454859.03100216,
  
    -39594.206766455, 
    -1830244.00548247,
  
    -58055.9638724756, 
    -1590154.142935,
  
    -182291.05050786, 
    -1592738.62950942,
  
    181894.429756595, 
    -1959341.81049234,
  
    321794.526287575, 
    -1410414.92446037,
  
    40952.696845411, 
    -3067228.3789562,
  
    251505.352277896, 
    -1750963.37391685,
  
    -91426.2611970182, 
    -3106780.14403558,
  
    -29376.7323713135, 
    -2851806.57238466,
  
    396337.250966195, 
    -1905084.16341996,
  
    -5594.575811715, 
    -1533792.49892462,
  
    33220.2285794095, 
    -1700993.65010145,
  
    483200.017436349, 
    -1904222.58699404,
  
    122328.828701501, 
    -1725333.88883745,
  
    181041.113019793, 
    -1780622.33763995,
  
    -161430.051673838, 
    -2268109.7399575,
  
    -156109.680492597, 
    -1750014.11393979,
  
    146740.308620572, 
    -2267870.49612625,
  
    265348.33566176, 
    -1035902.68148264,
  
    290086.469407607, 
    -2273184.38645492,
  
    244939.154504002, 
    -1302540.6841803,
  
    128390.222554609, 
    -1107775.66719881,
  
    85501.625688291, 
    -1615107.79111248,
  
    -250809.276208539, 
    -1261724.29195877,
  
    -28237.5923164864, 
    -2108625.27705632,
  
    -53310.5193606248, 
    -3074868.20073401,
  
    367871.756651591, 
    -1448081.43931493,
  
    -162085.810645429, 
    -1465161.91302769,
  
    333351.256149336, 
    -2488016.95359841,
  
    191572.670266769, 
    -1589071.93643677,
  
    166828.04497495, 
    -2440454.39645066,
  
    -275412.194432693, 
    -1465579.89768625,
  
    464003.801867008, 
    -1453961.27167438,
  
    20042.5960436057, 
    -2540426.61501299,
  
    40792.5094106127, 
    -2266866.80307087,
  
    326594.203630027, 
    -2212837.69935339,
  
    869.112148007293, 
    -2021786.75168189,
  
    398196.241296378, 
    -2369393.84991257,
  
    321299.869837088, 
    -2524620.38969256,
  
    366229.667180797, 
    -1146024.38689086,
  
    66477.0207009477, 
    -1015208.00573552,
  
    261851.374064444, 
    -1251445.54216663,
  
    431873.237229047, 
    -2266231.21086851,
  
    338406.921594665, 
    -2237144.23896993,
  
    -379616.583724739, 
    -1128812.4107427,
  
    -276750.849151663, 
    -1728535.61378398,
  
    292092.058047474, 
    -2582118.53711319,
  
    366971.41764342, 
    -1725304.56050527,
  
    217737.637498412, 
    -959050.842889122,
  
    465401.011047456, 
    -1653767.08003552,
  
    -195407.303755704, 
    -2704249.73293714,
  
    304012.692129761, 
    -2349893.10132767,
  
    -42919.811774966, 
    -3105898.59288975,
  
    507017.39733965, 
    -1455893.93787257,
  
    -217559.278789008, 
    -2735938.06391602,
  
    208051.084200108, 
    -2139013.98558483,
  
    312225.18250986, 
    -1293937.10390507,
  
    225171.891547471, 
    -1031948.30579849,
  
    278160.604844446, 
    -1920059.57224412,
  
    -214814.235427528, 
    -1091513.49797997,
  
    -226527.032733, 
    -1568467.7207826,
  
    126578.802321752, 
    -1327264.01636973,
  
    315249.934594158, 
    -1524044.88963945,
  
    80452.6871515029, 
    -2587893.61037138,
  
    -382182.409129419, 
    -1222581.14603772,
  
    276735.585829656, 
    -2197680.2317002,
  
    338222.883967725, 
    -1317160.02461721,
  
    332385.329656153, 
    -1067824.81715315,
  
    -65986.1089048168, 
    -2399648.31820561,
  
    -172236.312455259, 
    -2210113.89197404,
  
    303797.523314583, 
    -1113110.04752893,
  
    -19151.2924986908, 
    -3104836.55580439,
  
    -13738.6052293386, 
    -2941720.10803624,
  
    465464.216048978, 
    -2079112.89640504,
  
    -292977.154880382, 
    -1264404.68895133,
  
    98222.9879238301, 
    -1479188.05812795,
  
    -117866.477265549, 
    -2701772.89286557,
  
    307900.21565912, 
    -1250667.94624187,
  
    248786.544934547, 
    -1348675.65704126,
  
    197496.500907136, 
    -1777840.65723601,
  
    -67668.3443164803, 
    -1692575.69649927,
  
    -148439.116934416, 
    -1942282.68095108,
  
    -173509.373902285, 
    -2626482.25266363,
  
    157005.885678282, 
    -2574228.13262406,
  
    -47618.5118687172, 
    -2032402.37082325,
  
    117249.44827008, 
    -2065734.54168257,
  
    92251.2002607096, 
    -2669679.33393898,
  
    -264831.008270655, 
    -1675960.72742279,
  
    -245080.189358482, 
    -981933.311317329,
  
    -283537.354476796, 
    -1557124.30746248,
  
    113745.561877875, 
    -2778479.66295965,
  
    393452.592287481, 
    -1955151.9168583,
  
    -159778.293133659, 
    -2412945.74159035,
  
    -223231.019075507, 
    -1705084.72251964,
  
    -95231.4540199585, 
    -2937807.28318289,
  
    127646.076623966, 
    -2682892.53182718,
  
    295431.59238975, 
    -1240714.66369103,
  
    -88164.9009861152, 
    -1508417.09270909,
  
    199340.193582226, 
    -2356057.48006662,
  
    -69527.8533780157, 
    -1837996.20496686,
  
    137461.853070181, 
    -2083722.18737164,
  
    495602.33026799, 
    -2071242.88434936,
  
    -99227.9819057134, 
    -1355247.46180621,
  
    -180056.263034397, 
    -3052236.1994617,
  
    134845.156837378, 
    -2741914.6921094,
  
    178446.984414862, 
    -2111255.49569596,
  
    299164.812802678, 
    -1137371.79144127,
  
    -242990.971563756, 
    -1365880.49668316,
  
    76094.9581067569, 
    -2483866.72559448,
  
    252899.436883801, 
    -2117385.89026283,
  
    -73900.4240488929, 
    -2563264.7227735,
  
    -377485.561250948, 
    -1270681.25748628,
  
    -97704.7758604069, 
    -988359.823439481,
  
    -113900.635790059, 
    -1098852.26229694,
  
    270174.5727549, 
    -1500920.2825558,
  
    130248.697786329, 
    -1391263.75357547,
  
    257768.364959996, 
    -1718070.64057439,
  
    79094.0653466953, 
    -2105259.64782487,
  
    -246957.792095467, 
    -1598556.02983093,
  
    -101189.270828347, 
    -1690751.39706733,
  
    -100160.451691299, 
    -1317474.59901255,
  
    60766.0670891814, 
    -2876131.65702184,
  
    -72381.0850354094, 
    -2685260.33211106,
  
    7640.26380003756, 
    -2766665.94621121,
  
    -225010.402367529, 
    -1199850.95851704,
  
    -106698.909311078, 
    -2158596.08881995,
  
    217127.404012083, 
    -2656250.84390108,
  
    -62357.3831296212, 
    -1106425.22404813,
  
    481003.103986227, 
    -1602129.80537895,
  
    -293568.650216846, 
    -1381328.80077015,
  
    -41218.4138912161, 
    -1134833.96004279,
  
    -106282.307891548, 
    -1799032.40508558,
  
    292572.601335214, 
    -1889208.50736901,
  
    -344657.527646416, 
    -1379027.49251804,
  
    -220601.255723312, 
    -1148829.69346659,
  
    371376.196455885, 
    -2346008.20563792,
  
    36009.7271802116, 
    -1649234.63796586,
  
    113277.402107309, 
    -1395426.72504999,
  
    -164899.490812456, 
    -1241377.67819718,
  
    -106280.291007957, 
    -1081713.39223103,
  
    -18561.3234804353, 
    -2669279.98728014,
  
    161284.578334448, 
    -1365996.31255329,
  
    -126441.498371789, 
    -1266811.6008374,
  
    -120067.559692951, 
    -2785423.06614789,
  
    -217732.826142859, 
    -1458320.37799977,
  
    87906.6202386101, 
    -2000199.84081383,
  
    -66810.571692459, 
    -1005883.79641013,
  
    214196.886359823, 
    -2390722.86562572,
  
    449625.768776293, 
    -1480163.92197966,
  
    -127334.260681009, 
    -2053189.99022512,
  
    -94989.7907682705, 
    -2045952.87293751,
  
    -47138.0372447391, 
    -2172379.80727112,
  
    213128.903471985, 
    -1614202.5799138,
  
    -209427.229303403, 
    -1022242.11612192,
  
    53846.266623506, 
    -2775632.29795167,
  
    291257.663421766, 
    -1496444.57247091,
  
    24311.6424954687, 
    -2320558.67384772,
  
    -443368.928527814, 
    -1252674.25776488,
  
    253605.005621393, 
    -1488032.14716831,
  
    -122988.160470006, 
    -2154909.98935193,
  
    -160843.362732291, 
    -1552414.73222162,
  
    -398608.395300664, 
    -1296727.15905617,
  
    168279.570812455, 
    -1413046.71485568,
  
    -45920.7088743354, 
    -1533835.53368504,
  
    -60746.3710702894, 
    -1646581.87338393,
  
    359114.44041635, 
    -2352235.07855878,
  
    417985.434755206, 
    -2359559.57349087,
  
    -128558.790516035, 
    -2919826.16293676,
  
    -266437.203765358, 
    -1586123.04740629,
  
    -280495.796540617, 
    -1303383.68542196,
  
    24987.1449948346, 
    -1489902.18868827,
  
    -255895.087626448, 
    -1445940.51206092,
  
    400438.493515459, 
    -1872433.61606197,
  
    37442.006730043, 
    -1813434.98945741,
  
    -20307.7526602291, 
    -949379.618215054,
  
    468785.050785992, 
    -2233630.31132776,
  
    -11767.4542814511, 
    -2363837.3917947,
  
    175348.423962679, 
    -2618081.80237382,
  
    -170271.516366291, 
    -1796297.38867244,
  
    455401.584420851, 
    -2302652.89004269,
  
    350364.946322274, 
    -2366823.12111404,
  
    33018.7906318352, 
    -2451689.02176334,
  
    -52617.1786713393, 
    -2921177.69384506,
  
    81856.1704869126, 
    -1365670.39007433,
  
    418519.833508212, 
    -1072725.380517,
  
    -755.479343958497, 
    -2911286.04677498,
  
    174796.084452313, 
    -1651856.63535672,
  
    382900.338884581, 
    -1443238.84743495,
  
    -410574.428893949, 
    -1341684.92742157,
  
    92110.3255347893, 
    -2264141.6062056,
  
    248489.513940524, 
    -2390831.40645532,
  
    38580.8273217934, 
    -1992523.08481884,
  
    -204146.338134329, 
    -2005170.94650079,
  
    13055.2702841917, 
    -2264330.16489363,
  
    398501.793202224, 
    -2254460.37956962,
  
    629319.796667889, 
    -2204868.4886584,
  
    361395.367206785, 
    -1187713.45230074,
  
    -83970.7075148343, 
    -2301155.85833835,
  
    489712.221358757, 
    -1539110.81339887,
  
    244336.652576083, 
    -1551695.75578016,
  
    208782.370060026, 
    -1885721.22061317,
  
    -12007.5559305314, 
    -1574112.41948779,
  
    238976.684007847, 
    -1289095.92273107,
  
    131514.569050899, 
    -1215441.60267096,
  
    355644.43328011, 
    -1880209.25397521,
  
    -35255.7164897352, 
    -2242082.43453076,
  
    -251199.53758235, 
    -1715662.87115787,
  
    308199.179397343, 
    -1886290.47822521,
  
    -249658.577060248, 
    -1134349.21840892,
  
    593738.461122864, 
    -2224665.34230569,
  
    232709.744691916, 
    -2424089.69157634,
  
    166675.312943936, 
    -1464225.93999574,
  
    53495.7756367296, 
    -2535513.07607017,
  
    302674.809447126, 
    -1739592.52260724,
  
    338271.967975595, 
    -2373662.06707755,
  
    244975.110915313, 
    -2574885.04379976,
  
    330553.388468713, 
    -2030383.58698251,
  
    230583.857405905, 
    -2067351.88743314,
  
    283203.273692123, 
    -1389321.80808005,
  
    -75458.3498831392, 
    -1918078.75418534,
  
    189461.023824023, 
    -2153671.82336043,
  
    24517.0995426167, 
    -2363632.30274877,
  
    163506.11186461, 
    -928626.908225394,
  
    -476137.060259652, 
    -1332442.45920136,
  
    353011.500586075, 
    -1456620.78657748,
  
    329614.019017377, 
    -1502120.64906601,
  
    443899.74880455, 
    -2190825.80357172,
  
    80929.5656796349, 
    -2956350.71015312,
  
    -39799.2314675094, 
    -1935491.76034645,
  
    276020.24070287, 
    -2022131.9826993,
  
    120342.168816929, 
    -1898852.47700265,
  
    201320.329478516, 
    -2862792.57823261,
  
    -85615.1945549107, 
    -1561026.89311927,
  
    14825.2691561258, 
    -2083904.38559179,
  
    104035.82801952, 
    -1555369.15034109,
  
    -240421.797672872, 
    -1579925.94806715,
  
    390848.513034137, 
    -2016328.04364039,
  
    -60775.8310981145, 
    -2653434.24299291,
  
    124213.012119988, 
    -1570441.45192099,
  
    222203.487048227, 
    -1097340.03007128,
  
    -152011.392450562, 
    -2998974.26294467,
  
    63992.6676965575, 
    -2340689.49586383,
  
    -188741.099608932, 
    -1069914.15737383,
  
    135225.977924945, 
    -1261747.13375637,
  
    -3583.77123697812, 
    -2688689.09126289,
  
    375029.892234797, 
    -1306750.08884527,
  
    245587.313239387, 
    -2337310.10009636,
  
    297483.762681852, 
    -2101120.46895721,
  
    -30091.6814215965, 
    -1746027.60747489,
  
    99926.6980554844, 
    -2070864.44810736,
  
    356466.040480752, 
    -1937142.70906815,
  
    -302795.930625473, 
    -1622081.0620037,
  
    499207.787379709, 
    -2038739.73324643,
  
    -297225.304108313, 
    -1707205.65983619,
  
    334795.912097261, 
    -1137342.88001546,
  
    488344.294300411, 
    -2088923.15107642,
  
    24337.0162056246, 
    -1112773.64239332,
  
    -152883.364937335, 
    -1618015.6211444,
  
    269169.247684311, 
    -1296340.04645412,
  
    -29526.3538478231, 
    -2587594.96667436,
  
    121721.241003191, 
    -2167755.40089701,
  
    -146596.658084694, 
    -2662296.54812444,
  
    152777.6469216, 
    -2691661.00646811,
  
    167955.627619976, 
    -1894479.82437238,
  
    120167.873951537, 
    -2341288.05935657,
  
    244865.98973038, 
    -2187629.36281209,
  
    -62983.6859129634, 
    -1867237.01517897,
  
    -108588.419759368, 
    -2412774.02423143,
  
    -250732.106191544, 
    -1105891.02823909,
  
    18371.7338888082, 
    -1066506.57771501,
  
    -59506.6819465671, 
    -987731.148403518,
  
    -106231.503602677, 
    -2309162.08081517,
  
    136371.44184611, 
    -1419719.66401631,
  
    -16790.4018832466, 
    -2243801.70270484,
  
    -238204.387453592, 
    -1845062.89875224,
  
    149143.149136758, 
    -1839710.27246974,
  
    153503.371489184, 
    -1575099.51213211,
  
    218959.410835505, 
    -2303702.95579233,
  
    492318.526979126, 
    -1217754.05659697,
  
    28227.2464207715, 
    -2685673.22959054,
  
    -79972.6604739036, 
    -1063267.56241878,
  
    -22730.8530653655, 
    -1629891.29828585,
  
    116168.637314757, 
    -1993775.82190744,
  
    170364.547781674, 
    -2040904.57491373,
  
    -366478.825171957, 
    -1341896.6555788,
  
    435618.650037741, 
    -1899839.99096678,
  
    237206.699668138, 
    -1214764.16316559,
  
    505526.234496595, 
    -2016286.99724697,
  
    10727.6987849202, 
    -1529167.79172154,
  
    84587.5497686704, 
    -1299984.55040544,
  
    118354.819438198, 
    -1795018.95737428,
  
    -102001.778269839, 
    -1725734.72108288,
  
    126930.685662585, 
    -1976506.30010579,
  
    110911.638369988, 
    -2548643.96897226,
  
    109306.447093863, 
    -2715914.4371486,
  
    662713.887605077, 
    -2139293.26121369,
  
    13567.275058745, 
    -1626944.47590576,
  
    168061.040301945, 
    -1220202.53167414,
  
    -42254.1715759302, 
    -1411634.68248281,
  
    -32625.5208483524, 
    -1045471.60056294,
  
    190144.019745238, 
    -1071173.72101235,
  
    199410.7651937, 
    -1226932.90838336,
  
    -226860.35736817, 
    -1404996.70011402,
  
    14784.1923509152, 
    -3093687.57362904,
  
    310841.471626742, 
    -1354303.89867944,
  
    -121476.992573836, 
    -1410572.60664254,
  
    79398.3910662625, 
    -1098614.39352285,
  
    66291.557399207, 
    -2381809.44617997,
  
    -127843.856298336, 
    -1561467.04608064,
  
    62092.6145072418, 
    -1481786.20247653,
  
    115828.03792092, 
    -2873422.1054876,
  
    206412.264523264, 
    -1390120.75877797,
  
    -133737.840003815, 
    -1834963.1191802,
  
    -72718.1562129338, 
    -2509452.94293915,
  
    -55678.9945504349, 
    -2114540.25200128,
  
    178701.12895715, 
    -1168392.35716321,
  
    -19783.033474649, 
    -1435891.98827629,
  
    245445.615588079, 
    -1836095.34182885,
  
    -111584.182058682, 
    -1234419.21593005,
  
    -185540.955303458, 
    -2333560.54190809,
  
    235356.664153447, 
    -1861400.46725008,
  
    -73336.3789605604, 
    -1019123.00105657,
  
    -19218.8001549461, 
    -1713709.77955209,
  
    -131884.437403471, 
    -1375952.78734707,
  
    490828.993124409, 
    -1666380.3063572,
  
    25939.015503901, 
    -1914175.69628178,
  
    -79410.2150625674, 
    -1999112.02402315,
  
    231486.024302154, 
    -1633861.02345712,
  
    44384.8153096497, 
    -1593565.22377422,
  
    -22411.9397154082, 
    -2399988.89375762,
  
    294049.251459735, 
    -1572834.4657702,
  
    443102.555717497, 
    -1785221.93457179,
  
    37266.8232502269, 
    -2096498.8210709,
  
    -103921.996174468, 
    -1263347.65927841,
  
    76842.2322445191, 
    -2652871.66524688,
  
    225698.779118922, 
    -1734647.41887389,
  
    63583.4029537276, 
    -2095280.45515054,
  
    -264302.913149246, 
    -1812980.56660286,
  
    85553.0316499262, 
    -1704802.04568086,
  
    213123.362168837, 
    -1175104.3248058,
  
    -77130.1242270151, 
    -1465996.8178618,
  
    -40964.4562208799, 
    -1813640.15108173,
  
    -53000.9402885923, 
    -1608371.14793775,
  
    361769.411823984, 
    -1295380.61904588,
  
    250001.858187544, 
    -1767047.9660385,
  
    -199903.974909827, 
    -2913618.95472841,
  
    380591.447209179, 
    -1907106.1217158,
  
    372294.056862761, 
    -1792680.39376874,
  
    34101.20150627, 
    -1717329.14721519,
  
    483266.000907631, 
    -1890070.11247743,
  
    124812.038295152, 
    -1742240.93168719,
  
    178704.379373961, 
    -1763641.06523991,
  
    49868.1147517573, 
    -2941515.59118361,
  
    -146555.312148913, 
    -2260131.32223637,
  
    -156614.658484379, 
    -1766086.24503461,
  
    274449.477924726, 
    -1020977.70938109,
  
    378732.058163296, 
    -2427614.3560345,
  
    125257.296206642, 
    -1125138.54676334,
  
    81615.4057751387, 
    -1597531.09555498,
  
    -267207.533679627, 
    -1255629.23443475,
  
    -29602.1495919501, 
    -2092141.61057542,
  
    -58344.5031982843, 
    -3092229.45837007,
  
    383918.973206543, 
    -1457822.3089802,
  
    -25295.2985592176, 
    -2355822.44380084,
  
    -169744.812434889, 
    -1450766.2813559,
  
    189977.577356005, 
    -1569201.52767368,
  
    170967.689407637, 
    -2423716.88720993,
  
    -287057.222307792, 
    -1454281.93633005,
  
    7119.20016829556, 
    -2551895.00731247,
  
    328273.212765661, 
    -2196650.2122853,
  
    -301372.092129874, 
    -1691674.98863629,
  
    -6185.13793557012, 
    -2007112.53717917,
  
    405019.901654304, 
    -2384938.30758493,
  
    353904.527741633, 
    -1158407.94488068,
  
    258739.022739136, 
    -1267959.76052989,
  
    -270740.273084839, 
    -1167999.09758411,
  
    364845.640739102, 
    -1909128.07781463,
  
    -388381.664938012, 
    -1113888.93317717,
  
    396013.218710277, 
    -1235401.73624283,
  
    279894.756233626, 
    -2576113.50782889,
  
    -58548.846737528, 
    -2984633.9590611,
  
    234599.467152186, 
    -1950866.24415112,
  
    -207468.335354672, 
    -2690201.53216806,
  
    310718.454441989, 
    -2364965.53496043,
  
    -41134.2363739711, 
    -3122029.14273424,
  
    229962.197625248, 
    -2571041.64732269,
  
    361752.697103204, 
    -2004806.31402935,
  
    210478.44266329, 
    -2121741.57437634,
  
    307616.787872856, 
    -1310017.03011984,
  
    218853.760330129, 
    -1049339.91775871,
  
    582546.02470456, 
    -1575508.84513629,
  
    -199912.955324794, 
    -1098027.52725238,
  
    -220698.434010668, 
    -1585431.70037826,
  
    130457.914374816, 
    -1310659.23990799,
  
    311705.175233262, 
    -1506241.07067114,
  
    88589.3727372979, 
    -2573813.86621163,
  
    312143.27687219, 
    -2070308.65943708,
  
    -401718.525392589, 
    -1218462.14434653,
  
    276568.160723792, 
    -2214488.50681722,
  
    333136.735594784, 
    -1333681.85238452,
  
    319459.877471299, 
    -1079645.45594536,
  
    -75257.2038352631, 
    -2417498.04145359,
  
    -158309.6725739, 
    -2197330.15968974,
  
    -100531.947459822, 
    -2244392.60784743,
  
    321151.565854299, 
    -1103228.47448031,
  
    -20147.5846102631, 
    -3123496.59781828,
  
    -186715.17425171, 
    -2804621.77610086,
  
    107424.33890883, 
    -1496719.45841707,
  
    186130.585324197, 
    -2228925.86102967,
  
    182536.553555351, 
    -2256149.29189414,
  
    52090.8602860343, 
    -2377415.28492175,
  
    244271.873806032, 
    -1365653.6792053,
  
    121982.106397576, 
    -1018121.10005564,
  
    -53728.6539563988, 
    -1833398.01737566,
  
    -154094.306181247, 
    -1926550.57835961,
  
    -187335.226339921, 
    -2636332.35203182,
  
    154573.264078182, 
    -2590426.38237503,
  
    115253.613240255, 
    -2082375.74198219,
  
    -274664.115426027, 
    -1690452.36992385,
  
    100885.169140991, 
    -2886130.87024708,
  
    -288702.401349171, 
    -1541535.53481404,
  
    432722.314298214, 
    -1992909.73695541,
  
    111008.102434554, 
    -2793272.37537524,
  
    397894.690539459, 
    -1969078.3208546,
  
    83332.1100338947, 
    -2862343.54238856,
  
    -151195.556411262, 
    -2394920.31940392,
  
    -235178.304789285, 
    -1717804.51728798,
  
    193380.547474172, 
    -2373278.61890757,
  
    -69483.3944464565, 
    -1822178.33315873,
  
    137180.898120571, 
    -2101801.91281035,
  
    484829.250209549, 
    -2058270.16483298,
  
    -88757.6057271748, 
    -1369221.96237175,
  
    -165827.945475617, 
    -3057690.429294,
  
    147732.373724909, 
    -2749727.86096131,
  
    180790.080684588, 
    -2093143.78653015,
  
    315580.346693423, 
    -1127484.65168874,
  
    254236.830985818, 
    -2099264.88930981,
  
    -72146.227694151, 
    -2547503.41587759,
  
    -435464.46476946, 
    -1290713.77553622,
  
    -96987.636061137, 
    -1095323.92217575,
  
    369319.957110395, 
    -1974475.41312041,
  
    271372.572032645, 
    -1519004.77624182,
  
    135052.305283832, 
    -1374973.75809677,
  
    81096.8185476629, 
    -2088560.75762646,
  
    -215106.754271437, 
    -1248391.50876809,
  
    -99500.3142949859, 
    -1707757.14476152,
  
    -308286.705858569, 
    -1406972.54612015,
  
    -236270.012042102, 
    -1231397.13108099,
  
    -110844.196438569, 
    -1304489.01248888,
  
    58351.1298184635, 
    -2859612.84681434,
  
    -68273.1875247415, 
    -2668891.65561367,
  
    7413.39635782569, 
    -2781666.83931085,
  
    -241330.036014051, 
    -1194588.07705681,
  
    -16013.5382765662, 
    -2734354.28706552,
  
    -261912.160688524, 
    -1862166.72747801,
  
    202934.005170532, 
    -2661526.30197826,
  
    -45533.7442948794, 
    -1100879.33084686,
  
    467180.219863851, 
    -1617226.22898652,
  
    -307715.854569928, 
    -1385103.61772158,
  
    -58492.5706874205, 
    -1139276.07708978,
  
    4310.16199485512, 
    -1768847.96924894,
  
    -153672.145444491, 
    -2116864.9395613,
  
    -107920.486277667, 
    -1783661.60441597,
  
    373532.106905837, 
    -1265675.49715658,
  
    -236201.595015412, 
    -1144202.18462807,
  
    32899.3648828427, 
    -1631325.67243204,
  
    108659.942444313, 
    -1411450.30121361,
  
    -175264.952050834, 
    -1227483.79890583,
  
    158129.331246078, 
    -1382848.81362271,
  
    -116169.910497141, 
    -1280633.34643986,
  
    -224974.97795711, 
    -1443079.0639369,
  
    100022.343772826, 
    -1997195.60913925,
  
    -2566.03157647193, 
    -1714069.7690128,
  
    209866.391555307, 
    -2407348.33423604,
  
    466392.330729908, 
    -1489943.32936529,
  
    54200.1003627354, 
    -1791476.07290656,
  
    215023.067500985, 
    -1633451.1765969,
  
    -168353.19202932, 
    -2066406.55824461,
  
    60339.1802020316, 
    -2790155.47209671,
  
    287919.941055596, 
    -1478119.81857339,
  
    29640.4238877888, 
    -2302239.90866862,
  
    493114.795506453, 
    -1777605.83385223,
  
    29965.1254470607, 
    -1426192.42942722,
  
    230702.026932961, 
    -1457377.3330677,
  
    -166408.912333233, 
    -1537081.31016646,
  
    -416975.994544993, 
    -1295660.71597316,
  
    -150508.747899183, 
    -2534287.7113029,
  
    -46362.8230093486, 
    -1550416.76556158,
  
    366430.293636069, 
    -2367610.94772286,
  
    -133182.695768458, 
    -2935838.81003963,
  
    467110.260264821, 
    -1895796.07657207,
  
    -293893.093075731, 
    -1297651.2918168,
  
    28095.8356070136, 
    -1506873.84569845,
  
    -262660.839542755, 
    -1429732.70313536,
  
    237804.660669701, 
    -1995610.85840863,
  
    -43110.2913721012, 
    -2790445.28137206,
  
    182030.909978816, 
    -2603977.50176945,
  
    -168186.528886596, 
    -1812055.35515863,
  
    184726.14151507, 
    -1409504.09622989,
  
    480171.892245275, 
    -1416204.07670253,
  
    342800.273842489, 
    -2351441.07395565,
  
    31735.3961224416, 
    -2470962.51399516,
  
    -39681.4361985104, 
    -2893227.8348655,
  
    78804.7983337992, 
    -1382581.2898588,
  
    -156920.530505629, 
    -1035617.55034815,
  
    77388.9140703478, 
    -1494825.77698668,
  
    -28592.6294468817, 
    -2616951.13002735,
  
    -394218.614419063, 
    -1345784.42195179,
  
    91379.2121280568, 
    -2244130.83845774,
  
    243925.66141416, 
    -2407559.75833712,
  
    37712.0783919921, 
    -1975084.54777894,
  
    -195368.156084175, 
    -1992155.22987222,
  
    7177.81960541188, 
    -2190915.38196165,
  
    148540.200618356, 
    -1789030.76082592,
  
    375959.288851785, 
    -1176376.04388001,
  
    -122585.064369318, 
    -2425124.89081321,
  
    -25449.731959249, 
    -2011874.02021464,
  
    492604.108050504, 
    -1568987.87343569,
  
    241733.423294908, 
    -1532283.92008761,
  
    213630.742969576, 
    -1901223.75425689,
  
    556.861042730486, 
    -1646228.93689533,
  
    478295.857046344, 
    -2003949.08760267,
  
    126794.495317643, 
    -1232513.00214687,
  
    95909.5032154977, 
    -993061.767671683,
  
    -39718.9074683321, 
    -2261914.43596781,
  
    -239484.091169165, 
    -1703149.86404182,
  
    151029.495016313, 
    -985987.36516825,
  
    575880.574337156, 
    -2218737.85616663,
  
    44260.96612348, 
    -2550001.75395854,
  
    300006.781196974, 
    -1755935.89371609,
  
    328287.851002513, 
    -2359827.79235849,
  
    329964.867239105, 
    -2047662.24599194,
  
    228915.245618472, 
    -2049666.97622771,
  
    -188375.851677675, 
    -2491301.88696245,
  
    -82921.7677392092, 
    -1904806.49757298,
  
    136705.02609799, 
    -1632572.31521529,
  
    187217.292397707, 
    -2170269.55122785,
  
    169353.999764674, 
    -2512876.26155856,
  
    341310.726124868, 
    -1429700.62374675,
  
    325761.802299076, 
    -1484216.14185399,
  
    458982.692054883, 
    -2184027.44475085,
  
    273386.254919983, 
    -2039202.25400843,
  
    122671.901919874, 
    -1914990.90799578,
  
    51636.8951876122, 
    -1553680.50303582,
  
    -91978.1943297387, 
    -1544583.45859617,
  
    12808.1394592008, 
    -2100723.12809821,
  
    -52588.0550248088, 
    -2955406.86218094,
  
    106207.005643903, 
    -1573778.08941064,
  
    -235369.486285673, 
    -1594815.90893817,
  
    402715.487296374, 
    -2029657.41288615,
  
    121629.401120569, 
    -1551307.59494596,
  
    228916.095731213, 
    -1077298.20149957,
  
    -135973.782252795, 
    -2988864.73491697,
  
    60743.0134025751, 
    -2359161.26608244,
  
    -176210.716919369, 
    -1082646.68112059,
  
    -195810.740920323, 
    -1597102.10102011,
  
    140071.597548025, 
    -1244567.91698602,
  
    249992.649318029, 
    -2320802.87326326,
  
    300206.461395951, 
    -2084309.27544264,
  
    -286853.164652439, 
    -1354717.958225,
  
    -31386.1318193238, 
    -1729321.18175743,
  
    97801.2879710297, 
    -2088586.03906039,
  
    486942.796290009, 
    -2026462.86259206,
  
    -286668.452681793, 
    -1695771.51665684,
  
    317566.731464081, 
    -1148321.3949068,
  
    6472.66215566178, 
    -1116500.45302752,
  
    142986.634145524, 
    -2513074.66274167,
  
    -145396.385770825, 
    -1632380.07989817,
  
    -67392.7545075701, 
    -3110672.02951039,
  
    266022.314764845, 
    -1313037.75827455,
  
    319376.795310457, 
    -2121252.20563852,
  
    385802.423422822, 
    -1075092.98598662,
  
    -151555.628918536, 
    -2680269.2021253,
  
    163258.129691362, 
    -2677952.39780736,
  
    -335755.119769244, 
    -1078959.74555627,
  
    169848.001470965, 
    -1909203.81829482,
  
    258262.423473254, 
    -944202.763097841,
  
    116595.25663093, 
    -2359857.96761832,
  
    245021.546394896, 
    -2204824.44471892,
  
    -235893.777240227, 
    -1110059.21505788,
  
    700.829576836595, 
    -1069005.17667499,
  
    -43016.5080830779, 
    -984291.016752945,
  
    140492.150796808, 
    -1402669.29715635,
  
    -13358.3735058226, 
    -2225347.44038725,
  
    -250220.780058797, 
    -1836177.0474757,
  
    152665.832609545, 
    -1556780.87172536,
  
    214740.041717569, 
    -2320232.99205057,
  
    67392.6845966214, 
    -1865411.59834306,
  
    -97562.1810448126, 
    -1066937.03653231,
  
    27452.764346353, 
    -2637909.47366113,
  
    -20692.4963414225, 
    -1647580.99875397,
  
    167646.866419191, 
    -2181607.23494062,
  
    -341252.794082477, 
    -1344235.57056567,
  
    240482.078193822, 
    -1197384.91134347,
  
    516279.320238155, 
    -2031316.52634283,
  
    3365.81310984146, 
    -1512282.25700762,
  
    -215138.110760642, 
    -3019687.51096494,
  
    88409.8942246551, 
    -1282917.4339627,
  
    102705.038694733, 
    -1707754.29216618,
  
    108823.844790202, 
    -2565713.30447042,
  
    -213097.943821801, 
    -1972299.28977748,
  
    463797.962057472, 
    -1338193.28003738,
  
    16619.131382292, 
    -1646676.27584371,
  
    172078.206473523, 
    -1203284.74473764,
  
    -31453.6558821425, 
    -1424645.9478986,
  
    -13951.7158600311, 
    -1043159.6343525,
  
    197829.940895644, 
    -1051609.22888874,
  
    203639.69537397, 
    -1209726.79050649,
  
    191936.075071565, 
    -2523888.7006438,
  
    -238302.151320548, 
    -1392288.63218785,
  
    315662.200238469, 
    -1338027.5699512,
  
    -110122.299963048, 
    -1423885.00571571,
  
    96773.3111633747, 
    -1095880.52480731,
  
    19450.910966439, 
    -1846719.60674181,
  
    73889.2368557482, 
    -2365716.19191331,
  
    -127883.470413747, 
    -1577322.93654948,
  
    113891.627283762, 
    -2889667.54181278,
  
    202157.207712334, 
    -1406717.96479748,
  
    -135673.759610305, 
    -1818838.42022006,
  
    173978.258954316, 
    -1184781.73589244,
  
    322411.627532035, 
    -1723393.75014203,
  
    249487.745600615, 
    -1851106.85393516,
  
    -121694.847009501, 
    -1220721.12802418,
  
    -349046.183365444, 
    -1581715.42796394,
  
    -77580.6325342357, 
    -1320505.24207788,
  
    -78658.3082157169, 
    -2212092.99597063,
  
    -168570.15432007, 
    -2326471.65376869,
  
    230453.328719084, 
    -1844053.68255404,
  
    -82666.1242257465, 
    -1033286.52270122,
  
    -122287.165937697, 
    -1390407.33205856,
  
    707320.313320653, 
    -2142299.44078574,
  
    39117.9712955745, 
    -1928253.70392553,
  
    -81844.8841608341, 
    -2014093.10555237,
  
    227417.673006336, 
    -1614518.89702435,
  
    40965.4649808922, 
    -1575657.03222168,
  
    -31199.5639742908, 
    -2415991.54259203,
  
    292412.676494528, 
    -1553245.46167845,
  
    29053.0863674722, 
    -2247446.91500635,
  
    438788.526277916, 
    -1768928.94341707,
  
    36818.9247938874, 
    -2080098.47007925,
  
    -92914.2500710428, 
    -1276936.29920767,
  
    73253.2146493377, 
    -2668481.88602214,
  
    223525.628623488, 
    -1717279.7860915,
  
    61457.5480641554, 
    -2113005.74905553,
  
    -251555.443928984, 
    -1822163.03736175,
  
    68807.7442706357, 
    -1704060.47497696,
  
    209920.233254832, 
    -1192100.21079673,
  
    -42334.705675304, 
    -1797036.29668095,
  
    -47835.0440314517, 
    -1626987.71440743,
  
    356342.009804097, 
    -1312218.09159132,
  
    56907.7159072497, 
    -3044364.2968906,
  
    240646.995693246, 
    -1717675.21468948,
  
    -257453.406282496, 
    -1285601.51855088,
  
    -27349.022485943, 
    -1374411.37009479,
  
    -192752.640495367, 
    -2927533.56068167,
  
    380082.789056189, 
    -1932429.44405766,
  
    375320.112764988, 
    -1809505.99408718,
  
    34982.1744331297, 
    -1733664.6443289,
  
    176367.645728125, 
    -1746659.79283984,
  
    30039.6753851023, 
    -2964432.48708335,
  
    -145975.519547068, 
    -2240147.31417682,
  
    -157108.981241354, 
    -1781819.17303378,
  
    370674.112845567, 
    -2414338.68580026,
  
    122124.369858672, 
    -1142501.42632787,
  
    77836.8400176327, 
    -1580441.30144556,
  
    -283605.793347706, 
    -1249534.17962378,
  
    -30966.7071254476, 
    -2075657.94163943,
  
    400312.860142669, 
    -1467773.61140233,
  
    -25356.3678382761, 
    -2301114.5024775,
  
    -177403.813966312, 
    -1436370.65213913,
  
    188402.675271944, 
    -1549582.68698868,
  
    175107.336037319, 
    -2406979.37525607,
  
    30815.853459768, 
    -2563606.78906444,
  
    329956.811281294, 
    -2180418.4677261,
  
    -291266.120530258, 
    -1680323.75682849,
  
    -13124.1792574572, 
    -1992677.97782179,
  
    341126.931579759, 
    -1171246.10015531,
  
    -201362.501969344, 
    -2858076.071827,
  
    255626.671671859, 
    -1284473.98134817,
  
    -253620.380285949, 
    -1173358.69027593,
  
    437697.320871055, 
    -2508185.6016341,
  
    409298.073266838, 
    -1250287.72415829,
  
    -58895.4597987837, 
    -3000089.27730392,
  
    241411.251061834, 
    -1963807.36970068,
  
    317424.219209229, 
    -2380037.96833509,
  
    -288007.989877898, 
    -1067622.88813242,
  
    218632.406676079, 
    -2583583.10669942,
  
    374082.898102193, 
    -2016864.84455606,
  
    212944.514836076, 
    -2104193.67896848,
  
    303008.395948907, 
    -1326096.9585316,
  
    212347.174244115, 
    -1067250.27578409,
  
    -367490.559285078, 
    -1240033.14192657,
  
    -185011.675480092, 
    -1104541.55406977,
  
    -214869.8350303, 
    -1602395.68242893,
  
    342523.560243262, 
    -1497984.80826169,
  
    308229.69202553, 
    -1488785.20530026,
  
    96726.0583231043, 
    -2559734.12205183,
  
    312611.687128097, 
    -2052659.60712445,
  
    328050.587479873, 
    -1350203.68260686,
  
    306119.832286453, 
    -1091845.24891775,
  
    -84528.2985076583, 
    -2435347.7671565,
  
    -98268.0629244751, 
    -2226649.74347433,
  
    337958.286641432, 
    -1093658.55186103,
  
    -176142.586261388, 
    -1895429.99838613,
  
    488030.941890442, 
    -2104999.12152307,
  
    -116896.22170373, 
    -2738362.42725871,
  
    175430.561621213, 
    -2270945.30945579,
  
    239757.20241948, 
    -1382631.69891432,
  
    193173.548090327, 
    -1745550.27659846,
  
    127673.234212541, 
    -998859.915566383,
  
    -53559.1745875405, 
    -1816465.06409621,
  
    -201551.79322162, 
    -2646460.81526975,
  
    -117746.075077108, 
    -1357599.73440392,
  
    152140.639506992, 
    -2606624.62747393,
  
    113257.777952397, 
    -2099016.93982674,
  
    -301425.182139374, 
    -1541528.9687292,
  
    445253.860418752, 
    -2005385.61855384,
  
    108270.643249269, 
    -2808065.09024581,
  
    81385.5934393646, 
    -2879707.4236169,
  
    -145982.231735898, 
    -2933041.8926285,
  
    -142612.819688847, 
    -2376894.89721741,
  
    -350089.954283839, 
    -1402427.47815721,
  
    -246928.470021687, 
    -1730314.44440101,
  
    122263.618970622, 
    -2638962.71747736,
  
    323825.694830018, 
    -1883373.03400405,
  
    187516.818429866, 
    -2390222.59506138,
  
    -69438.9333179042, 
    -1806360.45863752,
  
    136905.157071053, 
    -2119546.06754679,
  
    474056.170409126, 
    -2045297.44777159,
  
    -78287.227093606, 
    -1383196.46267926,
  
    160815.640346171, 
    -2757659.88849611,
  
    183141.031465909, 
    -2074971.37004832,
  
    331517.096629007, 
    -1117885.8843749,
  
    103647.505970052, 
    -2475181.96765105,
  
    255581.896844128, 
    -2081039.94885415,
  
    -80074.6363322195, 
    -1091795.58205456,
  
    272608.98389369, 
    -1537669.1276759,
  
    139855.912781332, 
    -1358683.76261806,
  
    83102.5200414789, 
    -2071837.3020187,
  
    -245986.726051551, 
    -1249967.00765105,
  
    -250989.13306804, 
    -1226327.66523495,
  
    55936.1925477397, 
    -2843094.03660677,
  
    7186.52891561441, 
    -2796667.73241043,
  
    -257649.672373633, 
    -1189325.1933996,
  
    1785.53783590222, 
    -2736829.78141372,
  
    -248033.18669993, 
    -1870545.55492969,
  
    -28710.1079151681, 
    -1095333.43790364,
  
    453202.115921197, 
    -1632492.17980187,
  
    -75766.7247705697, 
    -1143718.19633377,
  
    5432.26566360165, 
    -1785735.61115463,
  
    -144641.127733596, 
    -2090117.33791994,
  
    -94230.6750467949, 
    -2783729.68264073,
  
    29846.0851453534, 
    -1613745.37751389,
  
    104042.483039346, 
    -1427473.87983225,
  
    -182660.86331964, 
    -1242488.23078744,
  
    233424.801326034, 
    -964590.913948856,
  
    154974.081444645, 
    -1399701.31249512,
  
    -155566.662271799, 
    -2147537.7953259,
  
    -232217.129771356, 
    -1427837.74987402,
  
    54768.1541859795, 
    -3114290.20300868,
  
    -2015.57133620353, 
    -1697999.8993893,
  
    205535.896492759, 
    -2423973.80039125,
  
    483578.720211863, 
    -1499967.60984673,
  
    -122005.04080591, 
    -2083417.41591163,
  
    53389.6028413548, 
    -1774239.5041108,
  
    216964.462613617, 
    -1653179.7534139,
  
    66832.0937805434, 
    -2804678.64624168,
  
    321795.576064024, 
    -1654581.37184108,
  
    -63870.7071474778, 
    -2883247.8549795,
  
    478452.759857397, 
    -1771355.95309712,
  
    -414106.56869735, 
    -1241337.54160388,
  
    19854.4604961764, 
    -1412494.34152135,
  
    -171974.461934172, 
    -1521747.8881113,
  
    -143744.65517991, 
    -2516627.12943851,
  
    -20405.0143676043, 
    -1542038.8971605,
  
    373676.41317212, 
    -2382840.2531371,
  
    -305810.929257759, 
    -1143933.42891912,
  
    514504.705284242, 
    -1818355.0433381,
  
    264480.368691985, 
    -2271427.14925408,
  
    31204.5237641682, 
    -1523845.50296664,
  
    -269426.591459058, 
    -1413524.8942098,
  
    419872.846280727, 
    -1901861.94926262,
  
    192206.837849381, 
    -1473812.72428781,
  
    756819.524149279, 
    -2041872.01892498,
  
    188713.398449988, 
    -2589873.20090701,
  
    -166118.177553539, 
    -1827687.58218868,
  
    187962.986759251, 
    -1392329.3078555,
  
    582918.611178273, 
    -2113851.86730902,
  
    335208.409077001, 
    -2336003.73806815,
  
    75753.4261806839, 
    -1399492.18964326,
  
    -169450.913195181, 
    -1022885.0266014,
  
    80207.3845717579, 
    -1509960.48236578,
  
    462808.98681651, 
    -2468009.42716473,
  
    -390745.965036534, 
    -1332686.21366623,
  
    25721.544080639, 
    -1976321.58820609,
  
    431552.214280939, 
    -2346591.62367909,
  
    -1416.39927432429, 
    -2264027.94075441,
  
    146262.815612878, 
    -1773222.38418641,
  
    643953.592954779, 
    -2224255.59595345,
  
    390123.731539688, 
    -1165349.61255736,
  
    -25905.9415214532, 
    -1995830.09776655,
  
    479210.795080652, 
    -1586963.48022195,
  
    239186.263986703, 
    -1513290.16657075,
  
    215177.3849063, 
    -1928147.40594341,
  
    122074.421842417, 
    -1249584.40407781,
  
    -102672.80995482, 
    -2428943.41325887,
  
    108341.016725315, 
    -975431.473396487,
  
    -49360.7167616836, 
    -2300395.40862898,
  
    -227753.175235927, 
    -1690620.33317306,
  
    145103.791239425, 
    -1007041.85030837,
  
    292344.077199104, 
    -1722200.1042057,
  
    318096.455943137, 
    -2345706.30852842,
  
    303604.037416601, 
    -2501388.1779286,
  
    227246.633831034, 
    -2031982.06502223,
  
    -183757.937760055, 
    -2521457.00179673,
  
    137205.942362624, 
    -1651473.59716414,
  
    184973.563168381, 
    -2186867.27638214,
  
    51583.9094558937, 
    -2007451.56558209,
  
    -235912.249137413, 
    -2901723.13048806,
  
    321974.741864111, 
    -1466614.48628583,
  
    474065.637760243, 
    -2177229.08567194,
  
    506967.597230047, 
    -2350389.54951419,
  
    270752.27159212, 
    -2056272.52505948,
  
    261255.065187964, 
    -1831028.79056665,
  
    -98341.1916495385, 
    -1528140.02381503,
  
    10791.0124753367, 
    -2117541.87280156,
  
    108385.704106353, 
    -1592250.79118065,
  
    -230317.174898471, 
    -1609705.86980918,
  
    414582.459361605, 
    -2042986.78484494,
  
    119127.546605697, 
    -1532779.22546954,
  
    235422.928160499, 
    -1057870.75473619,
  
    -119920.735517757, 
    -2978745.47775478,
  
    -258599.492249971, 
    -1069731.93213865,
  
    144917.219626126, 
    -1227388.69995764,
  
    454052.290561817, 
    -2482195.55807162,
  
    254397.985396671, 
    -2304295.64643009,
  
    -300714.944588705, 
    -1347558.31110616,
  
    -32680.5824750843, 
    -1712614.75358492,
  
    95679.3760427137, 
    -2106278.47193026,
  
    175635.843322487, 
    -1007744.12091303,
  
    -392180.599467107, 
    -1456021.69127656,
  
    299746.154562997, 
    -1159676.74956297,
  
    -11391.694607363, 
    -1120227.26146473,
  
    532854.390138546, 
    -1630739.00854463,
  
    -137674.815534703, 
    -1647194.62235539,
  
    -44887.1334667745, 
    -2611027.26277603,
  
    317675.300553401, 
    -2138527.4017062,
  
    -156768.615498728, 
    -2699162.47681839,
  
    156333.871124666, 
    -2412731.945902,
  
    321882.269968185, 
    -1007292.36538045,
  
    113067.721888107, 
    -2378193.55141097,
  
    262455.237902723, 
    -1990108.7933413,
  
    -221055.446091919, 
    -1114227.39916362,
  
    -16970.0771901628, 
    -1071503.775893,
  
    -26526.3342195921, 
    -980850.88510238,
  
    144612.862460563, 
    -1385618.93249339,
  
    -17630.4138156614, 
    -2185989.28577087,
  
    -262237.17046701, 
    -1827291.1934861,
  
    137349.563436943, 
    -1877006.39030928,
  
    151839.676613349, 
    -1538711.1657514,
  
    -85610.2864857521, 
    -1725760.76889377,
  
    62054.7443544128, 
    -1904491.2287629,
  
    -129989.155305521, 
    -1059312.17419331,
  
    -225760.606051231, 
    -927407.275925669,
  
    -42274.8705680953, 
    -1582833.93391947,
  
    168175.7180207, 
    -2164388.09942364,
  
    -341192.638230302, 
    -1363315.33520312,
  
    -3996.07256523481, 
    -1495396.72229369,
  
    -94812.0014979808, 
    -2834602.31778385,
  
    92269.3687381255, 
    -1265684.52942808,
  
    417135.668617768, 
    -1816491.22223803,
  
    105379.345956697, 
    -1725387.50208826,
  
    106736.051468452, 
    -2582782.64242351,
  
    84859.7166435929, 
    -2705453.05469172,
  
    -224741.509202681, 
    -1961961.65601553,
  
    248281.510494368, 
    -1688775.71567146,
  
    472565.800729246, 
    -1246462.43466563,
  
    4722.08667326234, 
    -1040847.6684001,
  
    205262.681503927, 
    -1032689.20290797,
  
    523363.816023025, 
    -2250884.14397429,
  
    129759.258769565, 
    -2018695.14451099,
  
    -249743.945530955, 
    -1379580.56180667,
  
    20525.7183568312, 
    -3074418.60249009,
  
    320482.928850192, 
    -1321751.24122296,
  
    114148.231260487, 
    -1093146.65609178,
  
    81486.9138572728, 
    -2349622.93790462,
  
    -122357.238712397, 
    -1722160.02023927,
  
    -166035.968469716, 
    -2507406.42486167,
  
    -137609.676503734, 
    -1802713.72345687,
  
    -51489.5728842841, 
    -2079609.01734601,
  
    334983.605033972, 
    -1693397.12170969,
  
    253522.091393852, 
    -1866089.45801473,
  
    -131805.511702282, 
    -1207023.04257335,
  
    -88716.0554075355, 
    -1306860.53632126,
  
    -80163.6083188439, 
    -2228741.80836904,
  
    -151599.35333667, 
    -2319382.76562926,
  
    52716.0335705845, 
    -2610983.98891236,
  
    362291.938134512, 
    -1830258.34923339,
  
    -7814.23102550585, 
    -2596090.97469989,
  
    722239.1713933, 
    -2116958.84788372,
  
    -84363.657758319, 
    -2029591.69052913,
  
    495679.217736557, 
    -1610627.59671965,
  
    513166.39043327, 
    -1919995.9971056,
  
    -124978.041391375, 
    -3157736.46502201,
  
    37630.604730194, 
    -1558191.36100318,
  
    -39987.190946219, 
    -2431994.18922938,
  
    290803.337573492, 
    -1533982.47186869,
  
    26241.2184384312, 
    -2230111.1006409,
  
    36371.0265955805, 
    -2063698.12154258,
  
    -81906.5015125873, 
    -1290524.93887891,
  
    56899.8936022481, 
    -2708935.20149562,
  
    420294.657987354, 
    -1964351.58647628,
  
    59356.5677662805, 
    -2130523.65645043,
  
    -238807.972253696, 
    -1831345.50786258,
  
    71471.8585171275, 
    -1720734.67206335,
  
    -43704.9526747023, 
    -1780432.44202211,
  
    -42572.9443705651, 
    -1645950.96805847,
  
    -177066.992648652, 
    -1557650.89868028,
  
    350914.60532918, 
    -1329055.5643948,
  
    -104813.162638402, 
    -1004141.08272916,
  
    -274065.734876951, 
    -1287707.31185714,
  
    -17161.9171109088, 
    -1388168.19351718,
  
    -161911.113426015, 
    -2928562.45083118,
  
    395869.171640647, 
    -1929661.95762219,
  
    378299.626518162, 
    -1826072.81525378,
  
    35863.1471019556, 
    -1750000.13898756,
  
    174030.91234032, 
    -1729678.52289476,
  
    331269.84853883, 
    -2510880.55025797,
  
    -145416.925730364, 
    -2220894.02172652,
  
    -157597.453837002, 
    -1797365.93332797,
  
    149117.731779623, 
    -2304231.49128831,
  
    217860.935552221, 
    -1217991.84146433,
  
    362584.91642572, 
    -2401011.52419005,
  
    118991.443768733, 
    -1159864.30834743,
  
    74070.4682870091, 
    -1563406.66721135,
  
    42558.7283375701, 
    -1872897.47649508,
  
    -10550.9187219372, 
    -2128400.36280536,
  
    -54475.0680493003, 
    -3118468.08841642,
  
    416902.632967212, 
    -1477843.81951399,
  
    -185062.815755764, 
    -1421975.02046734,
  
    186851.489975774, 
    -1530259.25825596,
  
    417532.526960797, 
    -1429975.35166806,
  
    34433.6633384674, 
    -2352390.52936988,
  
    331681.303339526, 
    -2163792.45511592,
  
    -281160.15112763, 
    -1668972.52773374,
  
    -19964.4831286871, 
    -1978448.80873223,
  
    527811.930576095, 
    -1560492.05471354,
  
    290337.002732627, 
    -2526057.22380348,
  
    327974.549632337, 
    -1184460.8217232,
  
    -189624.084355559, 
    -2846899.46283503,
  
    467991.774570312, 
    -2248113.60764727,
  
    -236500.487745092, 
    -1178718.28051272,
  
    84725.1390263117, 
    -2994076.13034447,
  
    -172678.63068944, 
    -1154027.86746772,
  
    389028.435986741, 
    -1397746.45001307,
  
    -59242.0704050121, 
    -3015544.59528864,
  
    323975.019209213, 
    -2394762.09417578,
  
    207302.615726923, 
    -2596124.5660761,
  
    386413.099101169, 
    -2028923.37508274,
  
    215471.216716983, 
    -2086214.37339563,
  
    298400.001569929, 
    -1342176.88720139,
  
    205648.568657808, 
    -1085689.2015804,
  
    -151330.873794938, 
    -1106669.46273135,
  
    201117.238963969, 
    -1903152.04674385,
  
    339987.489653756, 
    -1479647.4246559,
  
    304810.858358023, 
    -1471613.86144679,
  
    313087.244688549, 
    -2034741.31978981,
  
    -384943.490347489, 
    -1202145.15478711,
  
    322964.436651898, 
    -1366725.51063221,
  
    292350.579154294, 
    -1104437.56207126,
  
    -122586.203745356, 
    -1933521.83157083,
  
    -46499.6286887879, 
    -1863135.84088268,
  
    -96098.4715228196, 
    -2209645.88287976,
  
    354230.393299204, 
    -1084393.04398489,
  
    499785.543412234, 
    -1948827.83345077,
  
    450755.779063276, 
    -1700299.35614496,
  
    235242.531290956, 
    -1399609.72107837,
  
    191012.071552901, 
    -1729405.08505213,
  
    133199.388683439, 
    -980157.06165304,
  
    -203248.621412728, 
    -2671888.74265961,
  
    -106381.507820137, 
    -1369760.14930654,
  
    149708.017648863, 
    -2622822.87476973,
  
    -294330.331933751, 
    -1719435.65763897,
  
    -308982.913602179, 
    -1557111.17503476,
  
    457785.403826215, 
    -2017861.49795524,
  
    163919.906587096, 
    -2786759.59990314,
  
    -134966.381045419, 
    -2879323.25733031,
  
    -134030.082966415, 
    -2358869.47503081,
  
    -258527.793430062, 
    -1742663.77601666,
  
    -74846.2070772133, 
    -2910881.11696983,
  
    5591.37047014645, 
    -1975811.68104264,
  
    284579.755192546, 
    -1275461.16953083,
  
    320115.2100676, 
    -1866823.34537391,
  
    -69394.4743863432, 
    -1790542.58682933,
  
    463283.090350653, 
    -2032324.72825512,
  
    -67816.8511730918, 
    -1397170.96078977,
  
    185491.982247227, 
    -2056798.95356642,
  
    346984.673235288, 
    -1108569.70125114,
  
    18729.2306487157, 
    -2467085.46228355,
  
    256926.960505442, 
    -2062815.01111148,
  
    -63161.6366033059, 
    -1088267.24193338,
  
    411394.111886366, 
    -1698108.53283522,
  
    273845.396012765, 
    -1556333.48156499,
  
    144659.520020795, 
    -1342393.76468433,
  
    263025.962268077, 
    -1764153.75659293,
  
    85108.2215352951, 
    -2055113.84641089,
  
    -132211.685417027, 
    -1278517.8443516,
  
    383221.675876282, 
    -2530320.08703585,
  
    19630.4853769661, 
    -2798080.25692108,
  
    7950.4951726926, 
    -2677184.95465571,
  
    -234154.212453304, 
    -1878924.38483638,
  
    -11886.4693384694, 
    -1089787.54224737,
  
    -93040.8815667829, 
    -1148160.31338078,
  
    6554.36687732197, 
    -1802623.25331833,
  
    -111255.620963317, 
    -1752368.51464839,
  
    292900.655173808, 
    -1856954.50585693,
  
    26843.1530628223, 
    -1596454.9676526,
  
    119855.044436513, 
    -1423215.95772708,
  
    -171860.347625911, 
    -1255499.49620321,
  
    -63882.3709052005, 
    -1037738.93898385,
  
    -35619.1578365973, 
    -2702721.64469604,
  
    151818.834356269, 
    -1416553.81356452,
  
    -239459.281585598, 
    -1412596.43581114,
  
    89684.934334553, 
    -1967421.06159534,
  
    336237.373374087, 
    -1235742.44613862,
  
    -129100.649583155, 
    -1131420.82301983,
  
    201205.403885241, 
    -2440599.26628837,
  
    511907.221330427, 
    -1499927.00486062,
  
    363427.731198225, 
    -2514233.58076156,
  
    52579.1028649475, 
    -1757002.93557304,
  
    50836.9755409543, 
    -1003199.31264222,
  
    -196459.209102291, 
    -2045675.33667878,
  
    319594.651649254, 
    -1632975.52198632,
  
    463790.722011344, 
    -1765106.07505506,
  
    9743.79580332979, 
    -1398796.25607049,
  
    253521.665369214, 
    -1522984.69523712,
  
    144492.604775838, 
    -2840766.68864488,
  
    -174166.810834563, 
    -2611316.23497324,
  
    350217.729919909, 
    -1965083.58697694,
  
    -26452.3536205423, 
    -1527552.13251324,
  
    380862.943289105, 
    -2397944.31755371,
  
    404853.675157207, 
    -2332221.32983408,
  
    -275162.286899744, 
    -1537177.92901801,
  
    505010.195911841, 
    -1830532.41571885,
  
    12523.4913919711, 
    -1491994.93360174,
  
    43372.245523161, 
    -1519918.37757341,
  
    -46178.9900506605, 
    -970697.391105901,
  
    183788.393585204, 
    -1460485.4105272,
  
    -19137.2390857425, 
    -1933810.09044407,
  
    195395.884466142, 
    -2575768.90030254,
  
    -164079.590246295, 
    -1843094.86058949,
  
    191199.832003429, 
    -1375154.51948109,
  
    -226249.235255629, 
    -1332343.39053437,
  
    327535.681887711, 
    -2320401.97253043,
  
    241457.916846586, 
    -2236070.42818607,
  
    -127662.069637432, 
    -1883355.79565053,
  
    72702.0540275662, 
    -1416403.08942772,
  
    -181981.29808172, 
    -1010152.50556772,
  
    174216.289389647, 
    -1611048.22784555,
  
    -159781.371297855, 
    -1195572.65346144,
  
    422975.413583327, 
    -2332488.80176091,
  
    143985.430607398, 
    -1757414.00754687,
  
    384527.922341849, 
    -1152056.26464379,
  
    236687.143983091, 
    -1494654.64336943,
  
    272434.430488564, 
    -977107.282978657,
  
    229728.554886275, 
    -1338166.74806082,
  
    117354.348109154, 
    -1266655.80355373,
  
    -54358.3857343484, 
    -2318240.33297873,
  
    -216022.259302686, 
    -1678090.80230428,
  
    138978.797150521, 
    -1028804.426607,
  
    -199642.534747734, 
    -1140393.55633213,
  
    -237141.739351872, 
    -1350748.38005447,
  
    170298.863596316, 
    -1516254.39210213,
  
    288963.473201056, 
    -2506584.22176438,
  
    433713.171136522, 
    -1314023.89746588,
  
    155018.349425353, 
    -1651978.7280169,
  
    189502.315473547, 
    -2037410.62544199,
  
    -208671.186190327, 
    -2925188.98870572,
  
    489148.583465603, 
    -2170430.72659301,
  
    -319813.859496554, 
    -1638214.28617745,
  
    -46936.398867633, 
    -1901397.49589549,
  
    268118.285809227, 
    -2073342.79636851,
  
    382868.35692064, 
    -1696291.73436788,
  
    102931.866895098, 
    -2941100.32141898,
  
    265253.152767596, 
    -1846596.82200124,
  
    -104704.191424361, 
    -1511696.58929191,
  
    8773.88277841457, 
    -2134360.61530786,
  
    110628.266455627, 
    -1611264.99232726,
  
    -426879.928921138, 
    -1189878.57926609,
  
    426449.433623812, 
    -2056316.15409061,
  
    -61367.3693518923, 
    -2702656.04352919,
  
    124380.839033127, 
    -1492138.11006659,
  
    241728.05234575, 
    -1039045.54896887,
  
    -183036.039263184, 
    -3035936.85960631,
  
    -242779.631632583, 
    -1074006.47873492,
  
    -201797.012690824, 
    -1563059.30973144,
  
    149762.839249199, 
    -1210209.4831873,
  
    222389.054087885, 
    -2266856.85251726,
  
    137451.304435008, 
    -2616765.14635284,
  
    -33975.0328728106, 
    -1695908.32786741,
  
    93614.4902443994, 
    -2123495.40822206,
  
    575958.885904461, 
    -1528761.57691683,
  
    544821.991014223, 
    -2058523.82902691,
  
    183921.534979544, 
    -989928.393166232,
  
    -365872.347446041, 
    -1473099.16838431,
  
    462412.816307554, 
    -2001909.11857012,
  
    313293.336668519, 
    -1170616.23192798,
  
    450079.959132263, 
    -2051104.26969382,
  
    -505071.376499406, 
    -1326727.24225084,
  
    238879.203317852, 
    -1925303.74495526,
  
    -65353.3163494635, 
    -3078112.14564102,
  
    162688.756240427, 
    -1979518.25716045,
  
    315973.805796341, 
    -2155802.59777382,
  
    393002.320966422, 
    -1053523.5906052,
  
    -139972.910174447, 
    -2699532.19498221,
  
    160544.210035479, 
    -2395092.96963174,
  
    109576.771375016, 
    -2396338.97768117,
  
    326219.849440494, 
    -1807875.69413199,
  
    -206217.117140604, 
    -1118395.58598243,
  
    -34640.9815021387, 
    -1074002.37485299,
  
    -186155.778195168, 
    -2352881.0359043,
  
    148733.571411254, 
    -1368568.56563343,
  
    -279721.772044296, 
    -1782052.06785101,
  
    -274253.558420199, 
    -1818405.33923846,
  
    143733.065525003, 
    -1893743.55913645,
  
    151032.603118947, 
    -1521058.84745141,
  
    -85732.2055669796, 
    -1708877.08374224,
  
    70158.8206375477, 
    -1921411.04590519,
  
    137740.348666506, 
    -2173495.18328737,
  
    585814.651477855, 
    -2171200.98258198,
  
    168704.569622207, 
    -2147168.9639066,
  
    151885.869228182, 
    -2177704.30403574,
  
    47830.2941915479, 
    -3131952.88977607,
  
    -98540.6269358978, 
    -2699760.05188426,
  
    402363.323437287, 
    -1326374.04355429,
  
    -112395.277710743, 
    -2834059.46243371,
  
    96194.7477107918, 
    -1248157.35489996,
  
    422091.53041143, 
    -1833461.41776702,
  
    108053.650763632, 
    -1743020.71226834,
  
    104648.25788867, 
    -2599851.9779215,
  
    -205070.800039745, 
    -1963858.56308,
  
    219531.838068026, 
    -1499751.00290101,
  
    568446.072495416, 
    -1409434.79150996,
  
    23395.8892065541, 
    -1038535.70244771,
  
    64439.7698054782, 
    -2203414.69103308,
  
    503977.723009596, 
    -2223207.28869752,
  
    18238.7118744579, 
    -3057312.25810176,
  
    325303.659916936, 
    -1305474.91223668,
  
    21634.8580250399, 
    -1816395.95749638,
  
    89084.5933138311, 
    -2333529.68363784,
  
    -123216.178830173, 
    -1738752.83162523,
  
    -155422.020422554, 
    -1518549.92041959,
  
    329062.599881217, 
    -1976069.97966743,
  
    -139545.595852187, 
    -1786589.02695169,
  
    -43579.5321911586, 
    -2118135.28110059,
  
    -141916.17665309, 
    -1193324.95466749,
  
    -99851.4785388637, 
    -1293215.82810961,
  
    -49018.8492693738, 
    -1022194.73410172,
  
    365350.307288275, 
    -1846200.50344472,
  
    1166.07251233154, 
    -2583668.8740938,
  
    86410.2176620613, 
    -2544630.01502166,
  
    219429.121420763, 
    -1576538.98457323,
  
    -48774.815205074, 
    -2447996.83806365,
  
    40993.2150258962, 
    -2144330.04929915,
  
    -70898.7556671854, 
    -1304113.57635315,
  
    63430.0853744455, 
    -2696152.03246691,
  
    57255.5847553472, 
    -2148041.56164828,
  
    -226060.503033434, 
    -1840527.97862144,
  
    74135.9727636181, 
    -1737408.86914972,
  
    -45075.2021291255, 
    -1763828.58762127,
  
    345487.203309283, 
    -1345893.03694024,
  
    -6974.81419089619, 
    -1401925.0171976,
  
    -154152.491665481, 
    -2912208.97096455,
  
    381240.064703543, 
    -1842422.35337509,
  
    36729.0481015635, 
    -1766056.13704125,
  
    62757.4624723423, 
    -2447998.38276391,
  
    132112.811109656, 
    -1791948.58553577,
  
    171694.178694479, 
    -1712697.25049464,
  
    -144880.570126872, 
    -2202407.20519753,
  
    148502.918957496, 
    -2322559.02651927,
  
    213800.59090056, 
    -1234303.43708771,
  
    -119270.824079366, 
    -2649149.75535033,
  
    115858.517420758, 
    -1177227.18791198,
  
    70415.4712480243, 
    -1546875.74713544,
  
    -11730.1076993921, 
    -2110351.55864476,
  
    433685.075827111, 
    -1488030.9827763,
  
    -27945.2426087452, 
    -2337541.0297833,
  
    -192721.817545213, 
    -1407579.38879553,
  
    185338.426111991, 
    -1511410.73054088,
  
    39481.202054651, 
    -2335358.07673039,
  
    333405.795655788, 
    -2147166.44496072,
  
    -360646.089653432, 
    -1449551.87242496,
  
    479816.06240429, 
    -2238257.11538005,
  
    -219380.594946203, 
    -1184077.87320455,
  
    369012.103976607, 
    -1877980.99682361,
  
    -59588.6834662644, 
    -3030999.91353133,
  
    499422.111436912, 
    -1631350.51917933,
  
    330463.736093791, 
    -2409346.67588385,
  
    195972.824777779, 
    -2608666.02545274,
  
    217997.91885592, 
    -2068235.07027774,
  
    293791.606932913, 
    -1358256.81341616,
  
    233745.018262692, 
    -999361.641679131,
  
    337493.928567421, 
    -1461617.38279063,
  
    353208.077253862, 
    -1694859.61498626,
  
    313562.802248994, 
    -2016823.03245512,
  
    317878.288536978, 
    -1383247.34085454,
  
    -132430.381741464, 
    -1919730.00008402,
  
    -184833.807378314, 
    -2210183.97923307,
  
    -113654.480102685, 
    -2207194.36736419,
  
    -511214.720139301, 
    -1359061.69061451,
  
    53602.3411554772, 
    -2321827.58858735,
  
    52138.6459746496, 
    -889706.430856498,
  
    -189891.94663417, 
    -2687174.92161234,
  
    -95016.940821195, 
    -1381920.56175413,
  
    109360.132103465, 
    -2131515.36360413,
  
    -316540.645064981, 
    -1572693.3813403,
  
    153429.414863303, 
    -2773595.08012805,
  
    99631.5614407932, 
    -2870038.40473212,
  
    -139774.535280975, 
    -2897012.20155775,
  
    -377193.731987378, 
    -1400724.7260001,
  
    -270127.114641442, 
    -1755013.10491923,
  
    -98615.5515607896, 
    -2898011.02449502,
  
    6163.46983817615, 
    -1990690.53812194,
  
    316404.725305175, 
    -1850273.65674373,
  
    -69350.0129997552, 
    -1774724.71476309,
  
    136361.419162663, 
    -2154536.19561044,
  
    -57346.4725395139, 
    -1411145.46109728,
  
    361993.212683395, 
    -1099530.0006886,
  
    258272.026363743, 
    -2044590.0706557,
  
    -46248.6368743958, 
    -1084738.9018122,
  
    275096.162869716, 
    -1575214.51727696,
  
    149463.127518288, 
    -1326103.76920562,
  
    87382.1226953641, 
    -2158288.22277632,
  
    -257896.389689131, 
    -1536004.09275996,
  
    235362.250511723, 
    -2303953.9418434,
  
    -142895.432361274, 
    -1265532.260541,
  
    39042.7182746362, 
    -2232296.36722927,
  
    4937.16949625861, 
    -1084241.64904613,
  
    424877.885108388, 
    -1663426.00193646,
  
    -110315.038363001, 
    -1152602.43042779,
  
    7676.46809104228, 
    -1819510.89548199,
  
    286313.542471504, 
    -1841271.79166207,
  
    99779.9401960268, 
    -2975501.80208847,
  
    196460.803680037, 
    -936901.763390759,
  
    -147027.761985163, 
    -1821938.70003721,
  
    23874.0772717459, 
    -1579359.50650012,
  
    -161059.834387204, 
    -1268510.76187702,
  
    -46078.674827568, 
    -1037192.20052454,
  
    204499.307802064, 
    -2002620.20335562,
  
    102447.02550247, 
    -1797822.20174014,
  
    70771.2140323904, 
    -3115386.11980725,
  
    -111725.729486015, 
    -1128686.95430422,
  
    196874.9088227, 
    -2457224.73244345,
  
    -115204.5798613, 
    -1848231.42797771,
  
    51745.7616984559, 
    -1739280.60407679,
  
    113116.83648789, 
    -2918761.43052761,
  
    253217.888153078, 
    -1207551.4802881,
  
    -197273.336123425, 
    -2064797.17051223,
  
    368324.569894506, 
    -1356282.60361925,
  
    769309.508052904, 
    -2085659.64407263,
  
    317424.730950317, 
    -1611674.0283522,
  
    213667.23790671, 
    -1461538.27307569,
  
    -373985.08128727, 
    -1257454.20730163,
  
    -366.869147546424, 
    -1385098.16816461,
  
    254390.422430393, 
    -1541117.90467483,
  
    152125.433628069, 
    -2852385.20413852,
  
    -186797.951937738, 
    -2620047.82975271,
  
    214919.62050596, 
    -1818352.96859642,
  
    124271.761719638, 
    -1847201.9091724,
  
    -32499.6901604191, 
    -1513065.37006296,
  
    707483.563253878, 
    -2082826.25661724,
  
    396654.923154287, 
    -2318123.51904378,
  
    565310.813627497, 
    -2133075.82613152,
  
    495524.680833531, 
    -1842698.25392612,
  
    -65075.7667522958, 
    -2838673.73222988,
  
    202078.370482304, 
    -2561664.59969801,
  
    -162041.003197083, 
    -1858502.13653525,
  
    194436.67698957, 
    -1357979.72865167,
  
    -213822.643003534, 
    -1343481.17493897,
  
    319742.020343632, 
    -2304554.30042613,
  
    -34501.3356327081, 
    -2734155.75534295,
  
    -167078.856637302, 
    -2527898.28090564,
  
    172964.232612188, 
    -1591361.72735097,
  
    -149594.268377911, 
    -1209329.47714184,
  
    230429.865362155, 
    -2457027.28427278,
  
    414398.610430672, 
    -2318385.98010072,
  
    4116.42268976022, 
    -2227666.14834346,
  
    141683.870735097, 
    -1741437.82706886,
  
    441774.424741394, 
    -2230073.29076964,
  
    662198.277765746, 
    -2180972.1646204,
  
    -98222.9534973783, 
    -2373911.72046244,
  
    -147237.826544823, 
    -3148371.5600962,
  
    112648.495143751, 
    -1283675.77255242,
  
    -59356.0547070054, 
    -2336085.2573284,
  
    -283574.635631263, 
    -1767209.90930317,
  
    -228104.345309437, 
    -1365068.86034525,
  
    173572.282354751, 
    -1534524.41685912,
  
    297520.135244664, 
    -2317195.17943382,
  
    274322.906530489, 
    -2511780.26585816,
  
    328234.020646545, 
    -2098478.97178053,
  
    446054.793016891, 
    -2318536.19091192,
  
    152148.496931015, 
    -1632952.91051435,
  
    491884.726344385, 
    -2155518.29468308,
  
    265484.300026332, 
    -2090413.06767748,
  
    107466.526451267, 
    -2956135.02242687,
  
    269243.025439501, 
    -1862132.86317224,
  
    46593.4783855159, 
    -1908933.37751534,
  
    112880.635549862, 
    -1630362.31990534,
  
    438285.782056055, 
    -2069611.12779939,
  
    -61510.7058520464, 
    -2735892.38737533,
  
    115336.068565101, 
    -1475447.5286594,
  
    247835.766398718, 
    -1020809.75150334,
  
    -167465.501192316, 
    -3043142.43183221,
  
    265383.214699895, 
    -2610391.93522206,
  
    -204790.1499326, 
    -1546037.91298859,
  
    154608.461327293, 
    -1193030.26615893,
  
    91549.6041880514, 
    -2140712.34205878,
  
    559247.617347848, 
    -1531781.83880682,
  
    139951.873149477, 
    -1078106.36527692,
  
    27553.9303120297, 
    -3006266.08675717,
  
    437039.564128443, 
    -2038215.68352515,
  
    -107309.446867312, 
    -2497453.2634953,
  
    99382.1571446442, 
    -2789313.59359802,
  
    -163975.673445028, 
    -1641580.65358913,
  
    321189.554998749, 
    -1223653.11976391,
  
    256581.516006424, 
    -1363130.89373583,
  
    155458.146855896, 
    -1962830.20502527,
  
    314272.31129731, 
    -2173077.79629641,
  
    377954.615522636, 
    -1057004.33258799,
  
    164754.549204329, 
    -2377453.99581643,
  
    249074.478599017, 
    -970111.041794935,
  
    525544.113266091, 
    -1582897.58956767,
  
    106085.818664935, 
    -2414484.40666434,
  
    410835.548244757, 
    -1295615.28292126,
  
    331768.748231443, 
    -1822782.91200992,
  
    -115022.658102899, 
    -2387698.89338432,
  
    -191378.785734262, 
    -1122563.7725432,
  
    -168832.985962265, 
    -2345365.43520636,
  
    -269645.690301822, 
    -1769488.50790385,
  
    -188970.535010197, 
    -1868790.56423537,
  
    149946.929964453, 
    -1910035.94018181,
  
    -443193.709966691, 
    -1209006.6975623,
  
    -85854.1246482058, 
    -1691993.39859067,
  
    626020.065153915, 
    -2168714.98431349,
  
    523000.820262928, 
    -1431335.19854138,
  
    152265.539788972, 
    -2161220.86404071,
  
    -384716.181788355, 
    -1423790.45876588,
  
    -96135.6449390251, 
    -2680603.05766382,
  
    396383.382120479, 
    -1341359.1098064,
  
    309106.897121356, 
    -1945445.16294841,
  
    100120.124228429, 
    -1230630.18062988,
  
    426997.706920589, 
    -1850261.48173973,
  
    221638.4760961, 
    -1517784.12736288,
  
    42069.6917398442, 
    -1036223.73649532,
  
    15387.1055746752, 
    -2861241.78952715,
  
    461369.303019719, 
    -1177927.30078522,
  
    330124.388528651, 
    -1289198.58350844,
  
    18796.9707320876, 
    -1799876.48811902,
  
    96682.272770398, 
    -2317436.42937099,
  
    -124075.121402973, 
    -1755345.6432692,
  
    -149922.233295487, 
    -1533475.70124835,
  
    525309.471158057, 
    -1895523.61616814,
  
    -197823.447625916, 
    -2521015.9500726,
  
    -141481.513003647, 
    -1770464.32773342,
  
    -430286.210876541, 
    -1352797.57131614,
  
    -45517.9756498624, 
    -2099471.3191032,
  
    261319.267916792, 
    -1895046.32675752,
  
    -152026.84134586, 
    -1179626.86921667,
  
    -93495.3488272879, 
    -1433770.96839001,
  
    368366.121325678, 
    -1861920.82071259,
  
    -60542.4076599881, 
    -2035606.91000907,
  
    76561.527956315, 
    -2561198.8335739,
  
    -59078.0035757494, 
    -2260851.12297061,
  
    215581.637196912, 
    -1558246.92899339,
  
    36686.9581069976, 
    -2734467.69886581,
  
    -59891.0098217782, 
    -1317702.2138274,
  
    426067.895996374, 
    -1947862.366189,
  
    75546.1363185264, 
    -1895719.80410964,
  
    -213313.031358147, 
    -1849710.44912226,
  
    76796.2713240018, 
    -1754059.18444599,
  
    -46490.9212322702, 
    -1746673.75480746,
  
    -59215.273717104, 
    -1536067.79800973,
  
    545857.385913276, 
    -1492146.99583413,
  
    340059.798834355, 
    -1362730.50974371,
  
    3212.28898715424, 
    -1415681.84333305,
  
    -368832.00026265, 
    -1368918.0001508,
  
    37583.5164734874, 
    -1781900.18242019,
  
    57769.4927326277, 
    -2463800.72255409,
  
    149562.232044633, 
    -1467966.46700925,
  
    -180234.044247366, 
    -2268397.77339996,
  
    147888.106135366, 
    -2340886.56175015,
  
    209740.244051903, 
    -1250615.03542415,
  
    -119673.048306452, 
    -2665655.24428312,
  
    266813.548601564, 
    -1218675.84835071,
  
    266145.717142929, 
    -1107748.13241232,
  
    112725.59107278, 
    -1194590.06747653,
  
    95552.83215485, 
    -1650232.34883076,
  
    26221.6708871963, 
    -1878039.85503168,
  
    -12909.2939637884, 
    -2092302.7566811,
  
    450817.394585073, 
    -1498430.52545643,
  
    -200380.819076624, 
    -1393183.75957876,
  
    -254950.717549063, 
    -1502657.41658501,
  
    433336.144049192, 
    -1444101.46847902,
  
    335130.287714012, 
    -2130540.43235043,
  
    525537.889913164, 
    -1542343.31316333,
  
    451364.453794752, 
    -1897818.03267093,
  
    -211168.896094427, 
    -1171907.4891918,
  
    317608.227013017, 
    -1915193.95296014,
  
    -328487.187094479, 
    -1215261.32032593,
  
    336952.453236389, 
    -2423931.26004688,
  
    -29907.0189002886, 
    -3019432.16894758,
  
    205230.849021549, 
    -2070433.69829596,
  
    9026.36243692648, 
    -2421283.32516929,
  
    365946.280644163, 
    -1655827.14914679,
  
    282347.422404767, 
    -2162927.90051219,
  
    263470.482268433, 
    -1130849.10682931,
  
    365645.24954952, 
    -1024354.21814584,
  
    -38536.6731572003, 
    -1891719.07028742,
  
    -116619.37912975, 
    -2224659.98552044,
  
    -170596.704319592, 
    -1931527.90461424,
  
    485634.099123823, 
    -1934268.37919768,
  
    193005.173704074, 
    -2272129.98789276,
  
    54113.0788388953, 
    -2303044.15751103,
  
    -321308.284970314, 
    -1293332.71652117,
  
    87744.5963494587, 
    -1430083.24904633,
  
    542583.478225471, 
    -2242940.82421778,
  
    -176213.080204539, 
    -2702829.83350121,
  
    -83652.3711091899, 
    -1394080.97639872,
  
    107424.237730443, 
    -2147656.77105482,
  
    -282140.865048398, 
    -1710229.25139262,
  
    161217.116191239, 
    -2806114.53888657,
  
    -324098.376527782, 
    -1588275.58764582,
  
    142938.923139489, 
    -2760430.56035291,
  
    101598.768981856, 
    -2854311.53819358,
  
    -143937.465959609, 
    -2417667.78732342,
  
    312548.654622294, 
    -1833074.61563311,
  
    -46876.0963609577, 
    -1425119.96166281,
  
    -320360.578016523, 
    -1446647.03515428,
  
    185482.655354869, 
    -1906177.57015614,
  
    259617.092480073, 
    -2026365.13265489,
  
    -286980.199961873, 
    -1509004.31005281,
  
    404894.726314604, 
    -1732627.74449603,
  
    276387.947456197, 
    -1594714.74452966,
  
    154266.734757744, 
    -1309813.77127188,
  
    269063.002783767, 
    -1741811.5602581,
  
    -130417.583455274, 
    -2296715.16019325,
  
    229636.189362503, 
    -2320425.53228622,
  
    139518.520763415, 
    -1965250.66996342,
  
    48400.7961203734, 
    -2872769.33513686,
  
    371589.967849941, 
    -2541549.02582061,
  
    48025.7311688442, 
    -2199929.61067809,
  
    21760.8058759571, 
    -1078695.75610293,
  
    -161703.641462095, 
    -1130395.02720849,
  
    -127589.195159223, 
    -1157044.5474748,
  
    -118368.429404053, 
    -1959630.14620456,
  
    279712.005927297, 
    -1825554.73887432,
  
    -363978.719401901, 
    -1102028.88261865,
  
    54646.6931126448, 
    -1989718.08207573,
  
    -146329.912492917, 
    -1838146.12138459,
  
    20974.453591605, 
    -1562663.95162524,
  
    -150259.318435432, 
    -1281522.02974782,
  
    202585.930153794, 
    -991845.682268773,
  
    -75083.5543464811, 
    -1335920.32587863,
  
    102050.42407259, 
    -1780144.51573596,
  
    322753.575751487, 
    -1263190.15928679,
  
    -94350.809388879, 
    -1125953.08558861,
  
    -115611.361055156, 
    -1832598.79216679,
  
    -111498.040771601, 
    -1879328.5602956,
  
    248962.831342189, 
    -1224148.68630761,
  
    365177.636975045, 
    -1372980.31543966,
  
    742340.209462781, 
    -2096157.02351465,
  
    315300.236072804, 
    -1590818.45345928,
  
    200901.474226473, 
    -1456744.88105866,
  
    395760.691562, 
    -1178739.28388531,
  
    -10477.5338403851, 
    -1371400.08271375,
  
    -199861.869947147, 
    -2629078.59399093,
  
    232386.201948733, 
    -1897103.16595925,
  
    -8005.74451317569, 
    -1824213.92221762,
  
    -38547.0294133535, 
    -1498578.60541567,
  
    388444.109710463, 
    -2304004.96677288,
  
    486267.25413829, 
    -1854571.55087535,
  
    267342.942710387, 
    -1689840.18611561,
  
    44516.7524289064, 
    -1502860.59800897,
  
    -259317.579983788, 
    -992246.182527171,
  
    -63147.767930602, 
    -2854493.26224683,
  
    -446958.601120473, 
    -1388852.7367051,
  
    -276818.311676512, 
    -1802545.00470276,
  
    197673.522233742, 
    -1340804.94027726,
  
    -201396.050493401, 
    -1354618.9617986,
  
    -57800.0096985424, 
    -2569477.7614101,
  
    171742.616189755, 
    -1572153.89390587,
  
    -139407.163002935, 
    -1223086.3005642,
  
    225931.266850182, 
    -2473516.46122121,
  
    405821.809733023, 
    -2304283.15818243,
  
    139353.944098314, 
    -1725264.72842552,
  
    455797.168599077, 
    -2221649.81430222,
  
    -90102.2514240418, 
    -2356840.66466906,
  
    438390.27641549, 
    -1641750.04342489,
  
    1611.73042910514, 
    -1569726.4639522,
  
    223563.137108561, 
    -1370880.63144195,
  
    442373.512602281, 
    -1944216.77715912,
  
    108043.578384919, 
    -1300330.6822719,
  
    -46673.7027157096, 
    -2343599.27252599,
  
    -219066.951525029, 
    -1379389.33818101,
  
    304953.268522208, 
    -1413546.63787481,
  
    287019.23462371, 
    -2302644.83471203,
  
    259682.342314952, 
    -2516976.3096939,
  
    188585.996305788, 
    -2564844.3191714,
  
    448147.765217322, 
    -1325561.85835745,
  
    438071.771057937, 
    -2304641.99082522,
  
    70835.7097316623, 
    -1805818.15140969,
  
    476354.855593899, 
    -2163777.73338711,
  
    -54155.8826828359, 
    -1911387.02803488,
  
    273094.496724106, 
    -1877129.99191682,
  
    54638.3959665606, 
    -1924832.37491536,
  
    115199.476382903, 
    -1650023.26668542,
  
    449807.251681411, 
    -2082552.41619561,
  
    -37156.969232828, 
    -2661694.67265983,
  
    444066.364948237, 
    -1121932.48680941,
  
    253750.617664803, 
    -1003149.78362747,
  
    262467.26112703, 
    -2594168.08856423,
  
    -207783.286916338, 
    -1529016.51870074,
  
    159454.080950357, 
    -1175851.04938859,
  
    449931.195646445, 
    -2497560.03480686,
  
    332239.535724922, 
    -1380304.09135519,
  
    350567.140500794, 
    -1069827.8038327,
  
    423981.33113159, 
    -2025309.46750138,
  
    96306.6450414884, 
    -2772541.48893725,
  
    267988.236592751, 
    -1393941.07696839,
  
    253434.583086943, 
    -1379828.60555625,
  
    171187.686836431, 
    -2009627.10938796,
  
    312598.416759382, 
    -2190072.77617836,
  
    169086.634760537, 
    -2359304.98258561,
  
    538322.478988226, 
    -1573442.17346132,
  
    102594.86815185, 
    -2432629.83293438,
  
    337317.644567361, 
    -1837690.13014586,
  
    512257.917893315, 
    -2174467.16788748,
  
    -151510.193987379, 
    -2337849.83205337,
  
    -202870.451233078, 
    -1860323.26758803,
  
    -87552.9054805417, 
    -1873583.45168429,
  
    73858.3392887675, 
    -1910538.3060061,
  
    141585.688401041, 
    -2141432.90199817,
  
    415237.568180255, 
    -1996143.00472904,
  
    -111922.19121764, 
    -1019922.44670707,
  
    -93835.0290507982, 
    -2662277.4018909,
  
    390403.441061702, 
    -1356344.17851354,
  
    104045.503201089, 
    -1213103.00610177,
  
    431806.574714779, 
    -1866728.33609612,
  
    414865.759260886, 
    -1360503.784201,
  
    223776.724746912, 
    -1536087.84912425,
  
    434931.690852785, 
    -1265291.31558392,
  
    -80909.4312805271, 
    -3035440.23163135,
  
    -110417.209981712, 
    -2531264.0006882,
  
    -4006.7458618548, 
    -1434344.86002434,
  
    17423.1577256717, 
    -2843382.69955356,
  
    164637.391044676, 
    -2702343.11520304,
  
    334945.117140361, 
    -1272922.25478019,
  
    463839.247132832, 
    -1217703.44914226,
  
    -124929.394115472, 
    -1771848.27422556,
  
    -144422.446168416, 
    -1548401.48207709,
  
    -137102.39847407, 
    -1075097.81357595,
  
    514347.673990865, 
    -1889730.20142646,
  
    -143490.00850958, 
    -1753735.12484081,
  
    -71610.3396668291, 
    -1366422.59181945,
  
    -179795.906094125, 
    -1169814.25085233,
  
    189681.812723848, 
    -1214323.80926147,
  
    -75664.3227192692, 
    -2181011.67326563,
  
    43224.6414067772, 
    -2643645.39322797,
  
    -15371.5743130214, 
    -1011102.94550225,
  
    -21316.7676887638, 
    -1795370.85952846,
  
    -122208.017559591, 
    -1989558.84041169,
  
    -53716.9599044565, 
    -2240362.84022515,
  
    278717.654369142, 
    -1655048.57807574,
  
    437283.479585021, 
    -1960975.87448744,
  
    217020.981455364, 
    -1772276.8982781,
  
    79389.5654800096, 
    -1770290.13680058,
  
    -47911.10752089, 
    -1729464.77685412,
  
    -65420.4420034718, 
    -1520602.69829552,
  
    558238.740926955, 
    -1478892.69009295,
  
    201987.30363168, 
    -2232297.21497899,
  
    256136.777506449, 
    -1450505.31422456,
  
    13399.3943622004, 
    -1429438.66675543,
  
    387009.723308031, 
    -1874503.04119316,
  
    397128.351126778, 
    -1838640.52796159,
  
    52781.520795928, 
    -2479603.06505727,
  
    158293.839539751, 
    -1482975.41582066,
  
    479136.360722927, 
    -2219910.49008463,
  
    147273.295510226, 
    -2359214.0942679,
  
    205679.899400235, 
    -1266926.63104753,
  
    249246.676373681, 
    -1119363.33148096,
  
    -14088.4829412451, 
    -2074253.95252038,
  
    468027.632174172, 
    -1508877.36443027,
  
    282403.791340799, 
    -2494823.40622349,
  
    191992.281454425, 
    -2338709.77051129,
  
    232481.732582244, 
    -2664697.67828388,
  
    449174.888701568, 
    -1455315.39888201,
  
    336868.640945891, 
    -2113780.80845188,
  
    -358296.165205876, 
    -1433248.06379129,
  
    146337.493112254, 
    -2220796.13916737,
  
    144280.083712327, 
    -1180610.03133845,
  
    -226507.148476055, 
    -1170053.89315908,
  
    -185752.93628452, 
    -2295656.69267657,
  
    405640.895524912, 
    -1394344.79143638,
  
    -46724.3866399241, 
    -3014505.20897595,
  
    -104972.624004234, 
    -3187655.86793441,
  
    536759.430923442, 
    -1611641.30128221,
  
    395762.398536504, 
    -2467514.82802281,
  
    343351.293989431, 
    -2438313.82913037,
  
    -31317.6897039103, 
    -3000442.9091623,
  
    -387031.776206666, 
    -1241090.30580405,
  
    206115.884065782, 
    -2052747.67789088,
  
    -1238.32399701154, 
    -2439078.77067371,
  
    195684.279765183, 
    -1854456.3988837,
  
    364556.261913759, 
    -1634419.70698186,
  
    405655.601236092, 
    -1215590.35351082,
  
    283864.6301533, 
    -2145484.60474474,
  
    358484.464348438, 
    -1253586.4029994,
  
    373314.706190547, 
    -1040561.76753514,
  
    -119717.619836646, 
    -2242911.08930234,
  
    -164147.941875527, 
    -1947433.14895343,
  
    517039.614977271, 
    -1980510.44683233,
  
    199360.12159531, 
    -2258149.56202864,
  
    412248.743744926, 
    -1132992.88361443,
  
    92477.0261500802, 
    -1413305.32559641,
  
    109772.134785585, 
    -1008261.61688317,
  
    206822.178754904, 
    -2482566.8723248,
  
    312413.193857249, 
    -1979580.10918236,
  
    170590.950808673, 
    -2593788.11288822,
  
    97769.430945564, 
    -2652977.29458842,
  
    148023.834071621, 
    -2812304.95809496,
  
    480849.135656519, 
    -2075420.07979012,
  
    103565.976522921, 
    -2838584.67165498,
  
    270540.115285098, 
    -1327122.24135644,
  
    308683.056619524, 
    -1815833.08123883,
  
    -36405.7179854048, 
    -1439094.45951528,
  
    165611.910345848, 
    -2304480.78535255,
  
    -2185.70409348367, 
    -2953267.55491196,
  
    183645.35446973, 
    -1890827.83710492,
  
    243432.517943364, 
    -2029173.4878211,
  
    -55680.1235482733, 
    -2515355.57282578,
  
    -295889.751418903, 
    -1497145.72800937,
  
    277679.731784639, 
    -1614214.96932731,
  
    159070.339800203, 
    -1293523.77605121,
  
    271205.256995618, 
    -1722959.94439091,
  
    223910.128213286, 
    -2336897.12272897,
  
    170273.867274741, 
    -2225554.50953538,
  
    -144863.351955451, 
    -1161486.66452183,
  
    212793.134894611, 
    -914708.836378258,
  
    53701.0258129284, 
    -1972860.34248754,
  
    -145632.060545643, 
    -1854353.5424739,
  
    -139458.802999722, 
    -1294533.29270858,
  
    187844.285385825, 
    -2006123.96323959,
  
    101653.822900741, 
    -1762466.83218678,
  
    -117254.507493723, 
    -2940317.91268156,
  
    -116018.142249009, 
    -1816966.15635583,
  
    147807.499858837, 
    -2874481.03500138,
  
    244707.774789331, 
    -1240745.89478216,
  
    -180137.838977216, 
    -1993085.16331629,
  
    313218.321039639, 
    -1570380.86946691,
  
    420665.193055307, 
    -1734542.01726641,
  
    -20588.198791253, 
    -1357701.99480786,
  
    230713.707100288, 
    -1879880.55302779,
  
    340679.660351318, 
    -1939910.19524558,
  
    -9135.8820598514, 
    -1808546.19847271,
  
    477009.82744305, 
    -1866444.84782457,
  
    41506.7064970131, 
    -1486500.40025436,
  
    493257.667541823, 
    -1749126.30117377,
  
    213734.405871997, 
    -2534599.16669041,
  
    200910.367477909, 
    -1323630.15190285,
  
    -188969.458241298, 
    -1365756.74620321,
  
    -55913.9371907292, 
    -2554638.51672696,
  
    420594.501334834, 
    -2425458.11727558,
  
    170536.187919374, 
    -1553184.86493119,
  
    73196.1957693555, 
    -2786026.77776807,
  
    97267.8421686812, 
    -2210384.85225909,
  
    221432.668080178, 
    -2490005.63571455,
  
    -216282.823951517, 
    -1905198.30832069,
  
    137024.015006504, 
    -1709091.63004018,
  
    -65097.6072748535, 
    -1945423.6455643,
  
    423388.574269602, 
    -1395204.55111818,
  
    220480.425764674, 
    -1387237.57339055,
  
    103438.659429093, 
    -1316985.59470445,
  
    76328.7829255666, 
    -1647849.11883191,
  
    158424.482746688, 
    -1000631.59726304,
  
    86064.8259421886, 
    -3084256.09595449,
  
    56510.1623458779, 
    -2234608.25007578,
  
    70176.145331539, 
    -1789170.20089629,
  
    460824.984585381, 
    -2172037.16963611,
  
    300554.048148482, 
    -2541257.86495745,
  
    -66415.9795602886, 
    -1899832.68467638,
  
    -189256.874241827, 
    -2577608.5578409,
  
    57379.0797539298, 
    -1648158.51358327,
  
    276945.968008705, 
    -1892127.12066137,
  
    -46452.4286753671, 
    -3149793.26448642,
  
    -511301.420800449, 
    -1383459.69023217,
  
    461328.721306751, 
    -2095493.70459179,
  
    259551.307554155, 
    -2577944.24190633,
  
    -195320.052751515, 
    -1086830.11387175,
  
    164299.703286477, 
    -1158671.83481526,
  
    348700.558055867, 
    -1376684.79690175,
  
    308065.804134632, 
    -2223941.55331303,
  
    261747.753761955, 
    -1953747.61682863,
  
    -310123.57900827, 
    -1807839.59970164,
  
    534535.662365152, 
    -1478531.04756148,
  
    337231.130146804, 
    -1079593.57496869,
  
    410923.09813472, 
    -2012403.25147755,
  
    -89852.5418823368, 
    -2503502.69303347,
  
    93231.1329383236, 
    -2755769.3842764,
  
    -418234.559507283, 
    -1171748.26127504,
  
    272422.901565047, 
    -1378021.84098201,
  
    250287.650167458, 
    -1396526.31737667,
  
    310940.40327812, 
    -2206906.5320635,
  
    590393.271413537, 
    -2189712.90099284,
  
    173428.890137663, 
    -2341113.34685639,
  
    439526.771431332, 
    -1388332.8578507,
  
    342735.241854896, 
    -1852244.60986016,
  
    193796.223530741, 
    -2402283.63874358,
  
    427976.43335912, 
    -2008773.66864017,
  
    153024.883365571, 
    -2128253.98379245,
  
    -153806.260395322, 
    -994361.726436938,
  
    -91649.3754620406, 
    -2644867.489163,
  
    418462.253287678, 
    -1341420.6847007,
  
    125998.333179008, 
    -2565573.81477178,
  
    -86389.4474146541, 
    -3019492.07176429,
  
    -117420.121532251, 
    -2547045.10793539,
  
    -14690.4903511299, 
    -1421359.2759557,
  
    493915.340120039, 
    -1169290.31472844,
  
    -274933.438206508, 
    -1324440.36819044,
  
    -249531.762600361, 
    -1853047.22412007,
  
    172671.796139437, 
    -2690495.99682054,
  
    -125752.16170056, 
    -1787742.31261592,
  
    150363.900800911, 
    -1266728.62294774,
  
    -81975.8009052518, 
    -1352528.71252809,
  
    186526.563180479, 
    -1231176.31058892,
  
    -74120.4069932305, 
    -2165968.28775597,
  
    1452.06452167737, 
    -1005557.05230103,
  
    -21727.7729577748, 
    -1811368.82362712,
  
    213550.957771898, 
    -1954556.22516067,
  
    247592.349114364, 
    -2269845.54304738,
  
    -122139.073555143, 
    -2005037.59659784,
  
    -67629.5749385899, 
    -2001960.92309663,
  
    -48568.1987832285, 
    -2220685.8442191,
  
    207966.963897287, 
    -1522044.54949378,
  
    -7443.30245934291, 
    -1938517.69341104,
  
    -168388.392004972, 
    -1068385.02871231,
  
    13261.5840071592, 
    -2301956.92217074,
  
    445728.017279939, 
    -1834087.52989523,
  
    -37875.5178729153, 
    -1344879.49123092,
  
    275737.678580885, 
    -1635229.68281887,
  
    206404.259356737, 
    -1716884.36020659,
  
    87789.3731309593, 
    -1922627.23085214,
  
    81982.8620910417, 
    -1786521.08889711,
  
    193904.595533766, 
    -1277079.6350673,
  
    -49331.2965225681, 
    -1712255.79670376,
  
    -71625.610547871, 
    -1505137.59612627,
  
    -173045.431400977, 
    -1626008.05824837,
  
    -79856.3125745941, 
    -2736713.39234312,
  
    -262275.951787469, 
    -1297358.7998875,
  
    23586.4972822248, 
    -1443195.49043584,
  
    86198.9681352924, 
    -935057.910998102,
  
    394291.584618386, 
    -1821809.38677687,
  
    273347.258760481, 
    -2526082.82063857,
  
    146660.720880835, 
    -2377474.9074909,
  
    315602.307784146, 
    -1692317.7891586,
  
    485702.488468339, 
    -1519606.23263286,
  
    358836.701430305, 
    -2274685.12782582,
  
    -215698.822655502, 
    -1364392.49623515,
  
    266036.36096216, 
    -2497741.2584471,
  
    196267.262191743, 
    -2321425.07541515,
  
    246094.666430482, 
    -2652561.07274916,
  
    73870.4283329313, 
    -2262848.78537652,
  
    -12059.4987753859, 
    -2024993.00021751,
  
    39113.1460517701, 
    -911678.261236368,
  
    52016.4480755522, 
    -1839059.61891214,
  
    148168.815582331, 
    -1163710.82434398,
  
    -241845.403570744, 
    -1168200.29492938,
  
    -248503.881090057, 
    -1677230.08830045,
  
    -215449.93577343, 
    -1127457.11034976,
  
    30563.2576616999, 
    -2598753.07848881,
  
    406911.629767011, 
    -2476544.01619822,
  
    349622.962475268, 
    -2452410.55426175,
  
    178270.808157658, 
    -2645312.74978196,
  
    207000.916654985, 
    -2035061.65774378,
  
    -11503.0104309321, 
    -2456874.21617803,
  
    183050.752548597, 
    -1858926.56598585,
  
    363185.063792768, 
    -1613302.13742408,
  
    -195907.700442031, 
    -2402724.27694485,
  
    385647.855708718, 
    -1656375.79669956,
  
    -209983.875966438, 
    -2393803.41412888,
  
    -78920.4868648174, 
    -1647212.07918876,
  
    -122903.477910148, 
    -2261678.32080029,
  
    -240888.17239461, 
    -1535412.45434221,
  
    97209.4562087322, 
    -1396527.40460152,
  
    136361.611989869, 
    -943601.780645513,
  
    211070.362665438, 
    -2466648.51098047,
  
    178362.80248134, 
    -2578710.44316234,
  
    507911.582882026, 
    -2067765.01995441,
  
    469847.564695976, 
    -2062514.86035197,
  
    -119031.866250137, 
    -1035703.9183443,
  
    -355233.233188551, 
    -1417214.3631294,
  
    265860.236220292, 
    -1344342.59936397,
  
    -457664.13092772, 
    -1182260.29285438,
  
    -69212.4617683855, 
    -1725786.96771261,
  
    -529681.929811063, 
    -1214510.15557943,
  
    532594.617197885, 
    -2109398.28947155,
  
    -25935.3418068403, 
    -1453068.96008081,
  
    163129.716573755, 
    -2322740.37322931,
  
    181781.098358714, 
    -1875252.9098506,
  
    243594.945695746, 
    -2047128.30263431,
  
    323587.139642665, 
    -2276321.88445192,
  
    -304799.302875931, 
    -1485287.14596592,
  
    163873.947297686, 
    -1277233.7805725,
  
    279130.846785127, 
    -1757949.85640948,
  
    -259380.075437602, 
    -1569524.13319783,
  
    -89534.7439179802, 
    -1808098.37531793,
  
    218184.067064073, 
    -2353368.71317167,
  
    512325.072638886, 
    -1745088.22666636,
  
    -258940.840462452, 
    -930179.793579876,
  
    54008.7992887804, 
    -1436521.48388622,
  
    -132451.76271328, 
    -2833966.9324042,
  
    -4331.54489937746, 
    -2626367.27832025,
  
    182534.332553581, 
    -952436.787910558,
  
    67729.9797143771, 
    -2004033.47974906,
  
    -128658.289761, 
    -1307544.55838239,
  
    188486.25385478, 
    -1024772.6132567,
  
    47928.4369815518, 
    -2692563.68405983,
  
    -112633.979950891, 
    -2925316.60364177,
  
    -212314.533459983, 
    -1304073.41405719,
  
    -59600.9716496431, 
    -1120485.34841545,
  
    630740.05696558, 
    -2186261.7741822,
  
    139776.916349017, 
    -2583113.46628844,
  
    68496.767516716, 
    -1834953.53560867,
  
    135856.73969243, 
    -2884958.35011258,
  
    240452.717978435, 
    -1257343.10080168,
  
    -190262.631950425, 
    -2007160.01669117,
  
    479662.913511098, 
    -1702134.19939188,
  
    257044.374887797, 
    -1596512.77670052,
  
    376306.773658054, 
    -2503833.67317038,
  
    545983.99764057, 
    -1593539.49672767,
  
    273177.443604343, 
    -2243474.23364037,
  
    80853.8062451154, 
    -2206899.77410111,
  
    25061.6633827388, 
    -2137860.23181134,
  
    503129.056477421, 
    -1762988.73675249,
  
    452912.967762333, 
    -2401737.80051747,
  
    204147.212722074, 
    -1306455.36352843,
  
    -176542.865731158, 
    -1376894.53306284,
  
    -154266.317969346, 
    -2059869.33273362,
  
    -106878.365962467, 
    -1928373.80302241,
  
    -65993.1145189999, 
    -2597749.4238947,
  
    -159558.505392386, 
    -1050705.15764437,
  
    432440.26308876, 
    -2434945.41539856,
  
    73131.7899745107, 
    -2769439.25645868,
  
    -498496.743630854, 
    -1223541.75283743,
  
    453842.30521224, 
    -2366873.78815065,
  
    483842.651662433, 
    -2204802.86433841,
  
    -159984.348132839, 
    -1891406.51902342,
  
    217397.716875809, 
    -1403594.51508111,
  
    98833.7404732628, 
    -1333640.50713699,
  
    74662.2671658412, 
    -1627383.3582437,
  
    166542.528895464, 
    -984674.509907595,
  
    -35939.7817961658, 
    -2391973.94305076,
  
    428990.219973562, 
    -2458563.21371442,
  
    93949.2826444868, 
    -3100948.87514651,
  
    314944.369493762, 
    -2537406.91669082,
  
    -98594.0988757871, 
    -1565215.82731981,
  
    -189198.639414277, 
    -1649324.72274995,
  
    472850.190932074, 
    -2108434.99298792,
  
    -48874.7898590696, 
    -2689877.95066578,
  
    -134415.314487645, 
    -980750.232922444,
  
    -119762.257978957, 
    -3048935.49563393,
  
    274248.193841504, 
    -2601241.02091209,
  
    169145.322909533, 
    -1141492.61804494,
  
    324275.936840581, 
    -1433861.5612997,
  
    -356151.714031914, 
    -1320689.83710447,
  
    546836.489716443, 
    -1466525.51662644,
  
    -256355.011002128, 
    -1648268.62413056,
  
    397864.865137835, 
    -1999497.03545369,
  
    276857.566279305, 
    -1362102.6025406,
  
    280389.24115311, 
    -1229829.50951602,
  
    -57962.0780941777, 
    -1803773.32257154,
  
    571045.231657253, 
    -2190354.46199832,
  
    177771.147969817, 
    -2322921.71086907,
  
    -42328.6476073021, 
    -1982130.84495854,
  
    561678.026322693, 
    -1565669.33165402,
  
    121690.71304328, 
    -2809588.41617145,
  
    -203142.964413621, 
    -2742752.73428192,
  
    148848.620654782, 
    -1872939.51263882,
  
    189715.909769206, 
    -2418268.90556554,
  
    201817.655124496, 
    -2686608.80691531,
  
    440715.298537971, 
    -2021404.33255126,
  
    713041.529747508, 
    -2101516.31977633,
  
    153404.553668321, 
    -2111770.54134223,
  
    -142668.141472619, 
    -1005679.52411713,
  
    141337.339415456, 
    -1487556.76417113,
  
    133977.151767903, 
    -2548093.87984583,
  
    -92023.7722436102, 
    -3003094.84218841,
  
    -25374.2350984346, 
    -1408373.68943203,
  
    -127081.067871951, 
    -2523944.79740703,
  
    -289735.616963123, 
    -1318355.88333474,
  
    -264379.995503245, 
    -1846157.45195719,
  
    180706.201234207, 
    -2678648.878438,
  
    465782.346874398, 
    -1196649.66589047,
  
    10244.7764197504, 
    -1750093.80225758,
  
    89747.5501849548, 
    -2406766.60103445,
  
    -144216.303732856, 
    -1090883.57715429,
  
    -147527.918709373, 
    -1720102.45950568,
  
    -398619.684978308, 
    -1363245.72462039,
  
    145641.028343029, 
    -1283118.00193504,
  
    183371.3158341, 
    -1248028.80920331,
  
    -144393.173003081, 
    -1238637.00043113,
  
    -246122.60171638, 
    -1437339.79879353,
  
    208073.836338703, 
    -945266.986799153,
  
    33482.4641384491, 
    -992622.759556412,
  
    -22138.7782267852, 
    -1827366.78772574,
  
    -206068.428515202, 
    -1288978.44468565,
  
    215226.261094246, 
    -1969543.92142504,
  
    427320.056831831, 
    -1457459.68796866,
  
    -122070.132005719, 
    -2020516.35304199,
  
    204269.301276917, 
    -1504464.77039482,
  
    -179526.511185722, 
    -1057067.22857708,
  
    32206.0209059283, 
    -2780068.96940842,
  
    447910.736990694, 
    -1849880.52099317,
  
    48948.1791533001, 
    -2078001.8799103,
  
    208787.721379905, 
    -1735255.29019486,
  
    84576.1562470463, 
    -1802752.04125164,
  
    190701.466361708, 
    -1294075.51860323,
  
    -50751.4828111864, 
    -1695046.81875037,
  
    273171.566532699, 
    -1446344.37421657,
  
    400411.271431808, 
    -1097737.45180556,
  
    -163854.465504969, 
    -2871318.57676606,
  
    -413789.007440499, 
    -1380341.94806448,
  
    391415.972669783, 
    -1804747.7780211,
  
    431027.593868167, 
    -1699201.78641567,
  
    -185235.316261062, 
    -1683203.66989607,
  
    146069.147040511, 
    -2395109.70049595,
  
    -119621.270709487, 
    -2604643.97894758,
  
    320508.414113801, 
    -2331689.40589611,
  
    -75067.6760525086, 
    -2929525.53837622,
  
    -201076.072639674, 
    -1217295.40254546,
  
    249668.930325487, 
    -2500659.10821568,
  
    200542.242671029, 
    -2304140.37786391,
  
    488230.126659531, 
    -2189312.69017657,
  
    73879.0238965153, 
    -2242029.94428556,
  
    340408.594652722, 
    -2079651.74416416,
  
    4867.80106143261, 
    -2999238.33619183,
  
    27580.4055380549, 
    -918848.281387251,
  
    -24571.542224767, 
    -1500107.55179303,
  
    -145134.80775191, 
    -2740160.03577847,
  
    152057.547194297, 
    -1146811.61489448,
  
    347629.030424801, 
    -1818090.82360517,
  
    -188010.064618124, 
    -2314409.30626278,
  
    -258912.049349125, 
    -1691627.03058428,
  
    580021.73703388, 
    -1452876.17225102,
  
    355894.630703057, 
    -2466507.27693804,
  
    194558.166581877, 
    -2644335.09326848,
  
    -239792.103129311, 
    -1646332.57157771,
  
    1649.43648513656, 
    -2460794.87384505,
  
    361838.89232629, 
    -1592569.97383352,
  
    382309.314219425, 
    -1634854.56411889,
  
    559032.02736489, 
    -2246849.23379708,
  
    476691.706342816, 
    -1952864.10003571,
  
    101941.886009347, 
    -1379749.4811516,
  
    134204.91667698, 
    -925605.711225138,
  
    215318.546575975, 
    -2450730.14963607,
  
    272368.931050915, 
    -2550585.95438501,
  
    -107197.22956489, 
    -1606408.6515077,
  
    540165.951894878, 
    -1844833.5067926,
  
    136202.12698018, 
    -2047014.334949,
  
    -190236.119338293, 
    -1258149.97016964,
  
    243757.373448122, 
    -2065083.11744746,
  
    -87910.2905541423, 
    -1824454.63804464,
  
    214279.046759124, 
    -1336418.91881344,
  
    3739.03230735175, 
    -2323743.43507168,
  
    57831.1437447862, 
    -1419454.36744351,
  
    446105.860864327, 
    -1866665.84962945,
  
    -100010.155667354, 
    -1843873.22335507,
  
    -108900.487324253, 
    -3098111.28702449,
  
    -117857.774067248, 
    -1320555.82379818,
  
    181065.336999373, 
    -1042102.65425096,
  
    -44268.7885254571, 
    -1377385.55997297,
  
    -107933.56053427, 
    -2910055.91046523,
  
    -200959.840849232, 
    -1317385.81313036,
  
    -42226.049355525, 
    -1117751.4769868,
  
    132412.177202529, 
    -2596874.07751588,
  
    -114896.644536375, 
    -1569962.82637401,
  
    -200387.424665591, 
    -2021234.87252103,
  
    378329.244352179, 
    -1345059.19820298,
  
    -187097.625904215, 
    -1936505.5820346,
  
    -40809.5284349416, 
    -1330305.82145111,
  
    257950.76782265, 
    -1615431.54153644,
  
    505201.765189472, 
    -1856870.62925454,
  
    394830.201709919, 
    -2518962.26189647,
  
    324893.277508825, 
    -1942677.67922601,
  
    -11396.1568951692, 
    -1777210.75343783,
  
    -199065.345544904, 
    -1274770.97023069,
  
    27233.955352026, 
    -2119747.73966258,
  
    467482.627594148, 
    -2408596.9725974,
  
    207384.057708201, 
    -1289280.572699,
  
    -164116.273479048, 
    -1388032.31746745,
  
    -154232.452703881, 
    -2042966.49398466,
  
    -115928.976194874, 
    -1914755.15605089,
  
    -152097.98525873, 
    -1023860.26655655,
  
    -197248.859996126, 
    -2972058.91055124,
  
    444565.702751608, 
    -2444656.70806856,
  
    73067.384179665, 
    -2752851.73514923,
  
    248253.934924661, 
    -1093296.82088121,
  
    13182.0673128925, 
    -2701386.43913204,
  
    414549.411437414, 
    -2452515.49466554,
  
    94639.7207423489, 
    -3074709.43910062,
  
    55273.3246505367, 
    -2267164.36508045,
  
    448760.702844221, 
    -1165246.44799398,
  
    -146942.564265685, 
    -1582616.52041333,
  
    186059.903369523, 
    -2121815.03849376,
  
    -410385.689232476, 
    -1393581.22503972,
  
    331297.597940982, 
    -1557609.1267706,
  
    462765.927819322, 
    -1598029.70412159,
  
    -200526.640358754, 
    -2606415.98273146,
  
    -121243.481862608, 
    -1514976.08587472,
  
    -191008.121546409, 
    -1631724.11025644,
  
    -20799.6651773942, 
    -3066717.08183465,
  
    484371.658102353, 
    -2121376.28164203,
  
    -116757.349052188, 
    -3033752.818448,
  
    337708.015150778, 
    -1636842.26610838,
  
    277534.134149424, 
    -1950980.13310625,
  
    277764.220095881, 
    -2094412.36311272,
  
    330962.868341478, 
    -1024152.39768539,
  
    492944.938969181, 
    -1198202.45561402,
  
    174469.937717053, 
    -1027404.55250906,
  
    -118577.827046409, 
    -1142588.11867913,
  
    165078.931249553, 
    -2737331.02493585,
  
    -422509.363961425, 
    -1157223.39968981,
  
    281292.228796567, 
    -1346183.36681224,
  
    275874.570024624, 
    -1246807.53168007,
  
    349099.836982083, 
    -1911150.03611046,
  
    -149656.882528246, 
    -2624380.48251733,
  
    182113.405801973, 
    -2304730.07488166,
  
    -41940.4794217001, 
    -1998398.63997971,
  
    542216.150104026, 
    -2040172.6803372,
  
    101994.180369336, 
    -1047642.04418521,
  
    71965.5465966992, 
    -3090466.07853197,
  
    185635.596007673, 
    -2434254.17238743,
  
    147414.042842305, 
    -2092836.30624753,
  
    -98378.9075875193, 
    -2737536.15568669,
  
    132449.149206371, 
    -1471706.99919086,
  
    230448.879183461, 
    -1593202.43846912,
  
    -97845.9211374064, 
    -2986150.9950059,
  
    -36057.9820427277, 
    -1395388.10562142,
  
    -74700.2357798009, 
    -2999755.26230662,
  
    -76183.9535403171, 
    -2649156.62429098,
  
    -133964.571569885, 
    -2540665.72155578,
  
    -304537.795461703, 
    -1312271.40093407,
  
    194683.633087971, 
    -2698064.01203876,
  
    -103613.839785359, 
    -1108766.80477079,
  
    92908.9915617723, 
    -2389407.07623376,
  
    572751.278545566, 
    -2023953.42840519,
  
    -124358.980561048, 
    -2808729.96172348,
  
    -168931.562746384, 
    -2805902.10182204,
  
    -149546.872452736, 
    -1703286.12793657,
  
    -414688.770876469, 
    -1360264.90784234,
  
    140982.164221176, 
    -1299285.26018707,
  
    -155528.596134382, 
    -1224992.29221951,
  
    -236099.354582725, 
    -1450680.70247828,
  
    -195970.936588212, 
    -1302418.17047621,
  
    413114.149733111, 
    -1447299.74123354,
  
    -78866.7418698291, 
    -1952682.29344458,
  
    -4983.5210859025, 
    -1923059.99675773,
  
    -190664.630108433, 
    -1045749.43089688,
  
    50967.4511148912, 
    -2061165.26170215,
  
    211171.183661101, 
    -1753626.22263813,
  
    89352.8529692086, 
    -1906641.30393121,
  
    187498.33744768, 
    -1311071.40459418,
  
    -33383.9214015353, 
    -1546227.82916405,
  
    563073.092551322, 
    -1515571.30707358,
  
    -180702.583624993, 
    -2876160.70846864,
  
    388494.372513183, 
    -1787413.295356,
  
    74516.8902433157, 
    -2454965.58960884,
  
    432409.909797835, 
    -2241838.84161839,
  
    -131208.106501806, 
    -2204739.94061076,
  
    -183081.477695006, 
    -1699482.00480673,
  
    311809.607402107, 
    -2317357.89947994,
  
    -193945.557847278, 
    -1201513.69152792,
  
    400999.720893787, 
    -1436133.72420943,
  
    -113433.542841551, 
    -2128143.12783076,
  
    342178.572604627, 
    -2062587.2106637,
  
    211483.186123928, 
    -1849499.08052503,
  
    155946.27880626, 
    -1129912.40544499,
  
    342133.231493848, 
    -1802698.07694622,
  
    -170389.462501695, 
    -2307977.72454571,
  
    -269320.217608189, 
    -1706023.9728681,
  
    -266664.65142138, 
    -1118404.13276673,
  
    148130.0165722, 
    -2672818.6826078,
  
    -303953.316351376, 
    -1369104.87760672,
  
    69952.9977478963, 
    -2540071.54418939,
  
    210845.525006095, 
    -2643357.43675498,
  
    302624.344898985, 
    -1286273.07537867,
  
    360517.298044184, 
    -1572216.31840675,
  
    378094.30007791, 
    -1225073.18011508,
  
    379017.740172639, 
    -1613636.0918144,
  
    -398814.559289148, 
    -1144461.78797853,
  
    -87317.8562180344, 
    -1614492.89166718,
  
    -59125.5012568882, 
    -2184295.73747886,
  
    433351.47517524, 
    -1107248.08926455,
  
    106674.318523019, 
    -1362971.55989866,
  
    -68604.8154959197, 
    -2784352.81571849,
  
    -97811.299043152, 
    -971708.51202205,
  
    -140650.838515869, 
    -1614073.48349612,
  
    21507.6807849268, 
    -1783817.04145048,
  
    312950.825665817, 
    -2252260.62860838,
  
    -179312.922126393, 
    -1271205.81284798,
  
    90996.9179556451, 
    -1891040.05676537,
  
    -352661.783256408, 
    -1562495.23608783,
  
    446125.889507481, 
    -1281837.28567935,
  
    -86285.8396453287, 
    -1840810.90102935,
  
    217554.425284833, 
    -1319039.66699131,
  
    61653.4882007897, 
    -1402387.25100079,
  
    471333.435441113, 
    -2300154.36466019,
  
    -100290.719958736, 
    -1827230.83429433,
  
    362886.649018564, 
    -2317690.89613592,
  
    173480.743706141, 
    -1059814.93265924,
  
    -187494.916545857, 
    -2605230.10621005,
  
    174037.176230862, 
    -1330169.61150866,
  
    -189605.148238474, 
    -1330698.21220352,
  
    -24851.1292584018, 
    -1115017.60827122,
  
    125047.437798016, 
    -2610634.68628824,
  
    131878.863964965, 
    -2844501.13316667,
  
    383762.090127342, 
    -1330186.25363329,
  
    -179855.310419188, 
    -1952583.96527573,
  
    499616.287963757, 
    -1712877.87410234,
  
    -173088.459905291, 
    -2581585.66839661,
  
    364165.234596881, 
    -1210646.52705403,
  
    258878.984133325, 
    -1634805.83951833,
  
    516136.655723772, 
    -1847347.12612891,
  
    341593.277187584, 
    -1773244.59152243,
  
    -12526.2941838112, 
    -1761543.03214787,
  
    -189468.074079163, 
    -1289225.51494217,
  
    423759.612447188, 
    -2300955.64264601,
  
    295851.442964182, 
    -1634616.55499909,
  
    29030.1376924708, 
    -2932264.11491856,
  
    -45245.629415929, 
    -2837421.2977384,
  
    -151689.6809689, 
    -1399170.10432708,
  
    -154198.664396209, 
    -2026102.78691032,
  
    -13527.2172131139, 
    -1854930.02484687,
  
    695888.225559882, 
    -2174817.3075732,
  
    -474764.190175844, 
    -1215524.72498716,
  
    -143824.174374181, 
    -1887381.78378786,
  
    267881.201804974, 
    -1005836.71954546,
  
    256097.828841794, 
    -1075147.65286955,
  
    307241.147556296, 
    -1438022.49885264,
  
    -35752.9255557593, 
    -2323425.05349039,
  
    -36751.6145580513, 
    -2682873.82616665,
  
    -48504.3966453683, 
    -2407846.29475317,
  
    190893.47765918, 
    -1631199.7155199,
  
    182290.081469941, 
    -2352759.97041924,
  
    400486.277106009, 
    -2446625.93976648,
  
    464141.891182634, 
    -1157310.81473045,
  
    138575.902486779, 
    -1542972.80090506,
  
    333603.992429978, 
    -1576737.9486702,
  
    448355.429095275, 
    -1613702.1817283,
  
    349467.970535292, 
    -2551187.04261388,
  
    65839.041275128, 
    -1609618.34738836,
  
    -114801.568798583, 
    -1531908.68806033,
  
    464195.171336663, 
    -1430914.6687652,
  
    495893.12772764, 
    -2134317.57003807,
  
    221152.766876342, 
    -1999115.83335594,
  
    -113674.68016047, 
    -3018177.25806154,
  
    -256640.992844748, 
    -1042220.72409363,
  
    333804.370925925, 
    -1617235.91678626,
  
    262414.798632397, 
    -1922081.53079797,
  
    277588.744037862, 
    -2112028.83717306,
  
    -69856.6335564017, 
    -2439721.29257674,
  
    -5729.34324843337, 
    -3130981.52308331,
  
    -136442.183809461, 
    -1146314.92711639,
  
    285726.893768851, 
    -1330264.13082585,
  
    -41546.2920993718, 
    -2014918.60645744,
  
    396419.163871183, 
    -1284091.80516916,
  
    211146.95463156, 
    -1686255.10197834,
  
    -191690.735914014, 
    -2775911.55887336,
  
    173457.83325451, 
    -1266266.3710646,
  
    149402.609861052, 
    -2076255.7019773,
  
    -315848.905955262, 
    -1508693.97554864,
  
    -189533.658427686, 
    -1437031.983518,
  
    562188.551590797, 
    -1551702.14258508,
  
    250427.731159837, 
    -1948473.45148527,
  
    401656.994845803, 
    -1367797.34503026,
  
    151676.499014117, 
    -1726267.56390564,
  
    70982.0310620756, 
    -2138525.45305786,
  
    -245455.365660398, 
    -1881435.72126668,
  
    150522.190809019, 
    -895493.424201577,
  
    -122580.355096099, 
    -2576215.16283742,
  
    -121129.221870761, 
    -1113517.22537454,
  
    96070.4302255335, 
    -2372047.549236,
  
    -222073.435591523, 
    -1263840.84210943,
  
    -151565.828909156, 
    -1686469.79417044,
  
    -22768.3984963794, 
    -1057812.58015939,
  
    531783.005057065, 
    -1977945.04574903,
  
    177060.819202373, 
    -1281733.81160018,
  
    -166664.019265678, 
    -1211347.58400788,
  
    19562.8625881449, 
    -979190.998435809,
  
    -185873.442206192, 
    -1315857.89600874,
  
    -14322.2380762191, 
    -1891130.09324952,
  
    7102.54629178982, 
    -2357083.00536885,
  
    509263.411359506, 
    -1797360.57758971,
  
    -78354.529803022, 
    -1594396.29302435,
  
    406734.939665498, 
    -2436576.35843437,
  
    548274.562952972, 
    -1510486.30419543,
  
    534429.004810057, 
    -1945890.49378607,
  
    -11134.1578147199, 
    -2522917.64242762,
  
    -197550.701745001, 
    -2881002.8401712,
  
    -173654.516314833, 
    -2194156.27320029,
  
    154537.757463433, 
    -1712134.60799957,
  
    -180927.636673921, 
    -1715760.33945934,
  
    303021.476966141, 
    -2302879.22993175,
  
    -68340.7684101123, 
    -2950753.98864937,
  
    86462.5418962362, 
    -1559425.67930663,
  
    271846.863992366, 
    -2305217.3094012,
  
    462593.460455594, 
    -2207926.31708354,
  
    343976.113097375, 
    -2045256.93336711,
  
    -7915.29439126378, 
    -3000393.76436764,
  
    257936.331819914, 
    -1653106.30959819,
  
    295522.95432297, 
    -1820489.24633389,
  
    106075.547846066, 
    -3099338.22606196,
  
    60411.2482674159, 
    -2555600.29363722,
  
    312180.923527446, 
    -2512110.77458848,
  
    133877.483573277, 
    -1525879.51528983,
  
    368485.022474778, 
    -2224817.59625297,
  
    290018.577218878, 
    -2074732.82774125,
  
    -413263.584397062, 
    -1128978.76885681,
  
    -91396.8416847494, 
    -1598599.69301311,
  
    -16377.7199516355, 
    -2904342.09844514,
  
    -167637.331406076, 
    -2989274.72443969,
  
    -121530.093868376, 
    -3184175.01086717,
  
    -83129.7316935889, 
    -973479.347683884,
  
    20519.3250362179, 
    -1767450.91224368,
  
    23591.9197734772, 
    -2194382.20214738,
  
    -168389.724914489, 
    -1284261.65552632,
  
    -222383.292233939, 
    -1641912.79680809,
  
    -231125.96188399, 
    -1218856.0306529,
  
    290206.355816985, 
    -1442183.43666363,
  
    -258129.110624631, 
    -1618682.15716057,
  
    -139277.411370902, 
    -2151223.89233892,
  
    220829.806265564, 
    -1301660.41491115,
  
    -151146.096239897, 
    -2807177.07467523,
  
    -195879.251811223, 
    -2992029.81382498,
  
    65475.8326567905, 
    -1385320.13455806,
  
    433831.660989521, 
    -1838235.29889559,
  
    146388.724316499, 
    -2015177.96411651,
  
    -61417.3506595069, 
    -2218505.53890113,
  
    -185378.950965897, 
    -2104102.18408086,
  
    354491.522221156, 
    -2303493.7580851,
  
    511.990176041467, 
    -2841521.08289757,
  
    -178250.455627713, 
    -1344010.61127669,
  
    389194.936160533, 
    -1315313.31151862,
  
    219608.585039485, 
    -1865691.06074132,
  
    -179870.800158392, 
    -1303680.05939563,
  
    -73463.734144976, 
    -2038810.81427444,
  
    498833.697987286, 
    -1900828.04352165,
  
    -317828.664095303, 
    -1174496.83578049,
  
    -34456.9167956266, 
    -2452264.90684061,
  
    299239.832246136, 
    -1655068.53674562,
  
    31950.623822073, 
    -2918070.31183013,
  
    463746.189709857, 
    -1863187.70074725,
  
    462017.276227503, 
    -1752403.05710363,
  
    -139263.086261757, 
    -1410307.88847366,
  
    -154166.117057179, 
    -2009857.49050951,
  
    -34549.1028275393, 
    -2565136.60791396,
  
    -57489.5339524193, 
    -2424785.66209971,
  
    194572.185923947, 
    -1651731.80035065,
  
    19082.1283724288, 
    -2557807.53778381,
  
    64575.6564165381, 
    -2252092.32784224,
  
    370254.476694777, 
    -2305741.85492637,
  
    40322.7709291241, 
    -2798223.00721696,
  
    105780.384045802, 
    -1347917.63660405,
  
    335939.14691617, 
    -1596105.31022617,
  
    399089.847672269, 
    -2204870.51032125,
  
    61922.4888832638, 
    -1590668.70338088,
  
    -108359.653279529, 
    -1548841.28998789,
  
    450009.649500497, 
    -1421072.21036421,
  
    -110477.784677077, 
    -3002024.55199893,
  
    277415.88873563, 
    -2129382.29565681,
  
    114942.812340813, 
    -937672.109329725,
  
    -106579.344615115, 
    -2637590.39808549,
  
    290161.558483097, 
    -1314344.89238443,
  
    -62046.300059874, 
    -1756983.38190517,
  
    73158.0935293663, 
    -3149518.62829966,
  
    -186929.229508158, 
    -2368678.80114806,
  
    151391.179334824, 
    -2059675.09744899,
  
    161251.984887119, 
    -2501249.54321386,
  
    71134.6233722259, 
    -2154439.145738,
  
    -57425.4710212495, 
    -1369416.93748413,
  
    57537.1614620849, 
    -2652898.24606638,
  
    99231.8716023565, 
    -2354688.02443516,
  
    119358.754905285, 
    -2482877.24675525,
  
    340240.691364096, 
    -2278004.50241089,
  
    173905.571855984, 
    -1298586.31021457,
  
    -5279.73816042747, 
    -1793292.58210187,
  
    -175775.950279193, 
    -1329297.62179931,
  
    197722.693764246, 
    -1956949.01782651,
  
    -148827.37515132, 
    -1992305.72392605,
  
    -30848.7863438574, 
    -2176065.90428407,
  
    205816.661823303, 
    -1539895.14509634,
  
    5049.5338060169, 
    -2375458.36725306,
  
    65393.7542881985, 
    -2948941.2036413,
  
    181092.081816606, 
    -1345063.17386302,
  
    -65989.0075546157, 
    -1555721.82921141,
  
    570047.914348759, 
    -1483818.60624943,
  
    -93179.0795170328, 
    -2865222.76001582,
  
    -16444.4654815368, 
    -2539198.8306574,
  
    -423863.573880093, 
    -1370206.39364439,
  
    -178773.798107859, 
    -1732038.67436995,
  
    -133195.896103246, 
    -2682488.19770035,
  
    84744.1995831986, 
    -1542260.43216923,
  
    165685.486252618, 
    -1834504.496492,
  
    10477.7473380152, 
    -1918617.84774727,
  
    -405865.095251517, 
    -1323735.08349928,
  
    267175.393981995, 
    -2322340.12881216,
  
    -104309.589335047, 
    -2102100.76523576,
  
    345791.57500401, 
    -2027753.88414466,
  
    -430.565279387589, 
    -3016597.90110038,
  
    -233186.99817985, 
    -1128005.81332175,
  
    564160.605362031, 
    -2208131.01688996,
  
    243420.241854525, 
    -2641402.12372794,
  
    237180.258417058, 
    -2137264.35656907,
  
    198558.731594349, 
    -2086372.61746518,
  
    383567.968180126, 
    -2218019.23717414,
  
    69085.2948716281, 
    -2984575.74385744,
  
    585715.745474125, 
    -1492996.68835052,
  
    291577.015492142, 
    -2056815.5069374,
  
    80934.3000372927, 
    -2321799.92223898,
  
    -225260.572865515, 
    -1029103.85660282,
  
    -17710.3683512923, 
    -2704394.2647925,
  
    228063.098307603, 
    -2402975.0656025,
  
    15144.2743727147, 
    -2591200.44403646,
  
    -304521.158150155, 
    -1638910.96837467,
  
    473265.818513612, 
    -2021449.17152216,
  
    521581.020448006, 
    -2142147.69922218,
  
    -132681.207922224, 
    -2402159.02580789,
  
    -157466.527702579, 
    -1297317.49820467,
  
    103328.705819567, 
    -1919478.11472157,
  
    -188698.563892303, 
    -2190725.77266684,
  
    -25629.5894274947, 
    -1578499.25450991,
  
    224105.185049299, 
    -1284281.16554404,
  
    56893.4438630118, 
    -965556.920681793,
  
    69298.1746577634, 
    -1368253.01837337,
  
    70712.7019741372, 
    -1986912.03172253,
  
    433076.865685839, 
    -1347598.51892003,
  
    -181093.186726707, 
    -1455828.96987972,
  
    -1404.20843897785, 
    -2858044.36107133,
  
    -166895.763016947, 
    -1357323.01034986,
  
    462589.366023206, 
    -2394341.68202577,
  
    110352.889678749, 
    -2265388.05575769,
  
    355361.761537914, 
    -1404021.59064435,
  
    -14860.7405932968, 
    -1729179.32020394,
  
    -170273.528434607, 
    -1318134.60656214,
  
    430820.484015973, 
    -2318669.70572332,
  
    9884.69373117145, 
    -1883181.06100251,
  
    498872.627830564, 
    -1887172.58539579,
  
    124871.365892585, 
    -2711276.63798612,
  
    459739.978671899, 
    -1848057.2567207,
  
    445404.537701305, 
    -2415715.37727914,
  
    -126836.493751602, 
    -1421445.6753333,
  
    306992.732344952, 
    -2274757.91203857,
  
    -82430.0949789259, 
    -3098717.34547098,
  
    -180803.962744791, 
    -2930134.3856346,
  
    468637.333183546, 
    -1931755.13364058,
  
    134581.66811151, 
    -1775843.53452002,
  
    -77510.996404384, 
    -2837195.55116121,
  
    -523955.962372649, 
    -1195347.45209035,
  
    231814.520706869, 
    -1352859.58738404,
  
    -240477.110549344, 
    -1499473.78420988,
  
    377344.105218348, 
    -2321892.19407012,
  
    -207457.937585416, 
    -1634760.2008639,
  
    418708.075234366, 
    -1645945.86572445,
  
    58053.3803381833, 
    -1571948.60832257,
  
    200769.009068585, 
    -2190831.22166498,
  
    288112.008301817, 
    -1416678.35154728,
  
    350446.790353153, 
    -1283695.9020816,
  
    294596.223455373, 
    -1298425.65639804,
  
    -63451.8111885354, 
    -1740881.45993998,
  
    122076.078044737, 
    -2215310.94819172,
  
    86758.0246556398, 
    -3152960.87635335,
  
    -387549.479501693, 
    -1440337.67658214,
  
    121904.494025913, 
    -2749198.90140099,
  
    -197800.293606504, 
    -1679906.6666425,
  
    153379.746353569, 
    -2043094.49317866,
  
    -328982.902401177, 
    -1517246.20786429,
  
    285868.904887934, 
    -1740702.04156169,
  
    -494419.029468783, 
    -1345486.82300578,
  
    62047.0540234569, 
    -2639506.76446662,
  
    102393.310524156, 
    -2337328.49989228,
  
    339743.388857398, 
    -2303426.16031687,
  
    -56173.1538731613, 
    -1067372.90630622,
  
    170750.3223126, 
    -1315438.81154203,
  
    138890.141409263, 
    -2904085.74610057,
  
    -206029.615636764, 
    -1490703.41379056,
  
    73693.9727812809, 
    -1969646.98027895,
  
    -165678.458610222, 
    -1342737.34513485,
  
    199481.762129965, 
    -1972686.098917,
  
    -22493.4641452201, 
    -1901011.76538799,
  
    -163231.956397885, 
    -1587445.0481006,
  
    177888.955357594, 
    -1362059.05959593,
  
    -195500.599494954, 
    -1342658.58577355,
  
    557857.286360349, 
    -1491012.83638804,
  
    -302982.351230514, 
    -1513514.79551317,
  
    159561.741426965, 
    -1747769.31424931,
  
    -6196.87566629681, 
    -2303390.83292485,
  
    -176619.95708677, 
    -1748317.0090225,
  
    92807.3225649971, 
    -1505893.85836251,
  
    -387274.456146336, 
    -1319592.67006067,
  
    262503.923971625, 
    -2339462.94822306,
  
    -192622.185327864, 
    -1966164.7588369,
  
    -107825.161698568, 
    -2084977.98038313,
  
    347607.036910638, 
    -2010250.83492215,
  
    517908.722233234, 
    -1515685.65337267,
  
    -4750.84325375184, 
    -1628416.8928715,
  
    -285494.38910835, 
    -1752292.43796731,
  
    587279.001360351, 
    -2208973.28693134,
  
    -33524.2560631159, 
    -2515162.47372765,
  
    256024.477937897, 
    -2624039.61136085,
  
    235580.88964339, 
    -2120313.32403058,
  
    134791.556378852, 
    -1560370.62854491,
  
    196226.928409397, 
    -2103621.86230317,
  
    15677.2384755562, 
    -2446519.62094583,
  
    180318.027835816, 
    -934717.185146153,
  
    589192.948869109, 
    -1509369.00304522,
  
    293166.775119801, 
    -2038538.08066707,
  
    369492.479929692, 
    -1552233.41444107,
  
    -80576.1568596664, 
    -2113172.06796785,
  
    520547.573535318, 
    -2013757.31052736,
  
    86901.9188745269, 
    -2303360.71589873,
  
    232371.305261506, 
    -2386831.78305032,
  
    142100.908517628, 
    -2566861.52974194,
  
    -103103.276467117, 
    -1955778.45837116,
  
    18497.2905080604, 
    -1733968.14510712,
  
    -293960.987298719, 
    -1083499.55635083,
  
    -263136.231082893, 
    -1214987.65311545,
  
    -202155.216228958, 
    -1871720.46072097,
  
    532710.07726828, 
    -1458389.1714083,
  
    163952.752020422, 
    -2093020.49955671,
  
    -88646.9284482573, 
    -1052407.49842021,
  
    372195.214266429, 
    -1400884.08017098,
  
    -92203.1466366782, 
    -2177727.60931042,
  
    439397.284713589, 
    -2332772.52764154,
  
    -368278.681506434, 
    -1179745.69717526,
  
    -22600.4310523653, 
    -2439134.23460127,
  
    -185961.503081424, 
    -1858050.65647486,
  
    93071.3575632386, 
    -1752935.85985195,
  
    -158844.058292086, 
    -1011452.82606823,
  
    -187321.588348638, 
    -2245140.08638065,
  
    92550.4714215954, 
    -2593872.79550298,
  
    -252122.138424452, 
    -1488175.82285368,
  
    -319553.465848138, 
    -1542187.31780518,
  
    447676.635241729, 
    -1143084.1598353,
  
    384433.733741901, 
    -2338042.53321381,
  
    90257.5899257794, 
    -968672.208419073,
  
    -205874.639378935, 
    -1650160.73479317,
  
    403872.013242069, 
    -1662081.17692492,
  
    -190539.318577918, 
    -2749223.46561818,
  
    118820.578473649, 
    -1360473.57174825,
  
    -540515.178276571, 
    -1385401.53813215,
  
    182269.945231987, 
    -1829284.71472638,
  
    335788.541346964, 
    -1863390.12764763,
  
    543851.601458092, 
    -2022680.72726193,
  
    -86734.4842235504, 
    -2904444.12633447,
  
    107957.431159985, 
    -2674273.38621631,
  
    -75596.7329249246, 
    -1540325.62694642,
  
    -73547.3674311161, 
    -2091914.53293958,
  
    516906.930966642, 
    -2158339.99166342,
  
    -232440.858502112, 
    -1909218.85969344,
  
    230183.828319379, 
    -1687322.1685207,
  
    -106429.631288983, 
    -3042491.0326992,
  
    -217543.898606243, 
    -1876506.91419079,
  
    350442.700025668, 
    -2317828.88308656,
  
    -138280.091031908, 
    -2022183.3724846,
  
    -106136.994733261, 
    -2016591.80132961,
  
    59775.4527963708, 
    -2754263.38830824,
  
    174685.826443554, 
    -1379054.94558687,
  
    -207391.241926382, 
    -1330433.49403466,
  
    -70142.39354532, 
    -1611491.64579328,
  
    -242363.58379382, 
    -1478356.12991201,
  
    475227.789871671, 
    -2460969.94178752,
  
    162073.732181214, 
    -1765586.66750314,
  
    -174466.118520703, 
    -1764595.34393306,
  
    160719.430463113, 
    -2252423.79021903,
  
    60937.669250798, 
    -1498847.35031949,
  
    257832.453961256, 
    -2356585.76763388,
  
    -198856.504710439, 
    -1952755.28654489,
  
    465274.511951108, 
    -1471778.01906178,
  
    -7218.9115827295, 
    -1609947.48517228,
  
    -274062.772019031, 
    -1740082.58154584,
  
    252341.355597047, 
    -2607654.75550723,
  
    233921.080980751, 
    -2102721.70984381,
  
    -99426.1022337411, 
    -1909780.65659253,
  
    135259.780603307, 
    -1578038.282205,
  
    -60629.2232174798, 
    -2169174.04887008,
  
    75575.5290299257, 
    -1265332.79091851,
  
    155145.129140642, 
    -2144300.9341799,
  
    -160176.180664402, 
    -2653641.81773028,
  
    -232804.64477068, 
    -1097529.34543624,
  
    385270.902837134, 
    -2100397.21317354,
  
    -45147.5453485008, 
    -2992414.03980266,
  
    -113951.539192123, 
    -2042224.02467326,
  
    -178241.309432351, 
    -2013474.2734309,
  
    -2706.90468990255, 
    -1103143.99899397,
  
    -167561.516362575, 
    -3026256.64709353,
  
    -189405.331979728, 
    -1467453.78641138,
  
    -188382.307160897, 
    -1533892.90067897,
  
    341487.109441315, 
    -2470213.75515763,
  
    11922.1536924059, 
    -1349840.92520655,
  
    407716.627446023, 
    -2265074.61978702,
  
    -108039.229644217, 
    -1478075.85195903,
  
    367110.06698176, 
    -2167705.4763751,
  
    109970.993846855, 
    -1116297.16407253,
  
    -121027.864556155, 
    -2342362.40649335,
  
    475186.633565672, 
    -2145330.1566135,
  
    363482.196993176, 
    -1961769.78574797,
  
    340865.015531679, 
    -2388306.10760929,
  
    -100204.373412195, 
    -1166300.51833364,
  
    63872.9718335568, 
    -1323826.72269262,
  
    -267031.885976481, 
    -1553635.16921978,
  
    -102383.306624897, 
    -1138423.63519902,
  
    128845.866255952, 
    -1887929.43488349,
  
    100016.010467897, 
    -1622010.72236682,
  
    -56960.7737809681, 
    -1438745.58220452,
  
    32940.0793496459, 
    -1167152.36174044,
  
    109671.959137231, 
    -2212847.90280945,
  
    275945.402231977, 
    -2402440.69440367,
  
    217545.25344122, 
    -2432272.26152956,
  
    137873.367693627, 
    -2661785.93444926,
  
    228318.75607804, 
    -1966675.64556286,
  
    -97189.0524936403, 
    -1230717.45308074,
  
    134360.540497618, 
    -2425078.37831112,
  
    70879.8038954066, 
    -2707194.12822269,
  
    203788.715947524, 
    -2382000.7448507,
  
    -41281.3374264229, 
    -1262870.61269647,
  
    299919.218232858, 
    -2150643.60371431,
  
    69884.7221922903, 
    -1170104.70923372,
  
    221401.990009014, 
    -2146775.38062176,
  
    -51780.8026511926, 
    -1469112.72244223,
  
    92021.9229597846, 
    -1577109.69665561,
  
    -53177.8184568036, 
    -1948050.5262894,
  
    53577.4315143746, 
    -2801450.83054088,
  
    142168.250809448, 
    -1118844.03754941,
  
    47802.7302813751, 
    -1346545.88464918,
  
    385608.137099758, 
    -2196654.90194169,
  
    300190.541922574, 
    -2382736.33044921,
  
    487181.871350545, 
    -1826032.35273456,
  
    -178419.045383112, 
    -1397805.85435901,
  
    -213620.588222396, 
    -1399090.22984639,
  
    -297456.4763347, 
    -1572703.2307256,
  
    455505.4216654, 
    -1937985.95552887,
  
    -192874.924584691, 
    -1728480.13694073,
  
    -204786.23421527, 
    -1776855.78508246,
  
    103867.208513728, 
    -1079662.61765719,
  
    43576.1792126792, 
    -2706178.30090154,
  
    383236.624874006, 
    -1521330.50888031,
  
    331903.541330775, 
    -1053032.94405283,
  
    -134239.631325445, 
    -1704128.70404179,
  
    -208090.790293647, 
    -1755822.71844595,
  
    449848.458701821, 
    -2206237.80893699,
  
    -44289.9424819798, 
    -2524038.50707928,
  
    34465.6516566162, 
    -1376675.59462551,
  
    -265123.12851509, 
    -1782657.14210962,
  
    -77473.8744659657, 
    -1127844.65814811,
  
    -45838.324199232, 
    -1451774.50808936,
  
    -190749.781220874, 
    -1830882.903497,
  
    452640.111586071, 
    -1532214.1731773,
  
    -165237.255661825, 
    -1709523.23505449,
  
    -83053.1114622161, 
    -1201471.06415256,
  
    83636.0135888787, 
    -1127137.74082076,
  
    409609.940769104, 
    -1836050.97286431,
  
    45042.6729050214, 
    -1251882.27538907,
  
    49590.8934467786, 
    -1136149.76504524,
  
    531151.768412232, 
    -1597269.445812,
  
    -4662.63362609597, 
    -2545546.92156899,
  
    -312300.785029789, 
    -1664530.4271509,
  
    368206.481621608, 
    -2446650.28916674,
  
    443737.149485405, 
    -2115829.31718712,
  
    369299.649388778, 
    -2244286.93520954,
  
    278876.220887427, 
    -1046838.37884536,
  
    349768.684960067, 
    -2412471.393346,
  
    -198166.009570855, 
    -1818412.68487449,
  
    434330.448006893, 
    -1816761.72547147,
  
    402022.443931042, 
    -1530712.26003565,
  
    -4981.79341146768, 
    -1321642.6027395,
  
    -68169.1017074267, 
    -2015171.76017132,
  
    -173551.628297636, 
    -2398822.29940191,
  
    -185646.798509543, 
    -1790700.63942473,
  
    187694.917419128, 
    -2688356.44769343,
  
    98226.7352062897, 
    -1291624.05947383,
  
    39056.1663268417, 
    -1050115.85872367,
  
    385351.530276793, 
    -1476465.84118611,
  
    399747.685204843, 
    -2050319.77931865,
  
    -211247.723350746, 
    -1574245.50505486,
  
    66141.7354737818, 
    -1047587.18735136,
  
    -190329.380441218, 
    -1765410.8716707,
  
    583553.983624674, 
    -2241675.42097603,
  
    411919.742729448, 
    -2217819.70411776,
  
    21432.747594854, 
    -1370141.25718401,
  
    -86261.3528926857, 
    -1981924.2429605,
  
    -284142.167257413, 
    -1235483.93795067,
  
    -251060.060564175, 
    -1421164.56947325,
  
    475332.169954686, 
    -1546892.12111731,
  
    56851.5260205973, 
    -3094497.03051807,
  
    -160261.05846268, 
    -1411570.28856779,
  
    -135461.116529373, 
    -1687573.11425604,
  
    18336.6468372354, 
    -1301585.24845308,
  
    140211.860803308, 
    -2687276.7717317,
  
    -74312.1621057703, 
    -1260573.75256908,
  
    374824.930241159, 
    -2070317.50813477,
  
    14637.0928509386, 
    -1098507.64571972,
  
    340925.431744614, 
    -2212863.00998248,
  
    370674.354002953, 
    -2099057.58329046,
  
    -159584.237043843, 
    -1437280.15039516,
  
    275101.979535458, 
    -1987598.30399812,
  
    -54979.11482647, 
    -1992045.88564216,
  
    -140953.74857556, 
    -1674470.83712207,
  
    -229351.342208189, 
    -1734815.08746216,
  
    53351.1482718221, 
    -3062200.786567,
  
    -96525.3429159142, 
    -1787953.28194106,
  
    -163002.522060604, 
    -2900192.88592098,
  
    -71567.1497661196, 
    -1075767.40230509,
  
    -166638.966294287, 
    -2230914.76097566,
  
    359375.580023281, 
    -1011198.17512455,
  
    -200534.957768256, 
    -2804837.23944658,
  
    -290676.35737445, 
    -1610095.05821428,
  
    -58434.7619786294, 
    -1975640.3554166,
  
    72257.4662143544, 
    -1288840.9836585,
  
    135814.296377753, 
    -2331802.357908,
  
    543771.772379626, 
    -1448067.81612775,
  
    628341.476628979, 
    -2227319.53217247,
  
    288619.278846618, 
    -2352123.99263746,
  
    358121.773806, 
    -2039812.41738439,
  
    -255055.794564234, 
    -1703644.95222762,
  
    -79645.1533427692, 
    -3083371.79312895,
  
    -81445.7239583357, 
    -1426229.1351668,
  
    -107875.523226887, 
    -1217167.43753903,
  
    -415147.894036998, 
    -1274432.53847703,
  
    -93669.5311557422, 
    -3038965.6333928,
  
    443800.301528109, 
    -1588717.7801409,
  
    -220196.774498005, 
    -1430391.91514808,
  
    170286.008373717, 
    -2559595.4526922,
  
    43318.9292844404, 
    -1277213.24447429,
  
    -82935.5280488829, 
    -1245387.44848766,
  
    -175020.547762356, 
    -1850572.75988871,
  
    79652.2924549549, 
    -1188952.3691252,
  
    3625.60374115872, 
    -1152667.0315196,
  
    -408524.561724223, 
    -1158105.02611233,
  
    306330.735463952, 
    -2418542.23803325,
  
    369064.520508308, 
    -1466450.99677509,
  
    425242.864484379, 
    -1613680.15192902,
  
    90797.8254331664, 
    -2813633.45654373,
  
    411502.66736429, 
    -2372248.94434947,
  
    -151459.381046527, 
    -1334081.09406811,
  
    -141553.707803608, 
    -1508296.70082684,
  
    215468.001976199, 
    -2189763.93710339,
  
    260806.723357221, 
    -2175653.11984267,
  
    367895.134579734, 
    -2116829.57413601,
  
    293754.282129973, 
    -2210697.52066788,
  
    -388046.98073083, 
    -1283704.20852926,
  
    -144489.586461991, 
    -2068429.18001109,
  
    230270.700791489, 
    -2200160.03867097,
  
    -157683.720684402, 
    -2635802.43058983,
  
    -224196.599715292, 
    -1484529.77185128,
  
    385936.326135752, 
    -2376117.05288137,
  
    131007.139189403, 
    -1759218.664348,
  
    237328.44256505, 
    -2603811.36148523,
  
    259091.023195928, 
    -1554014.62002911,
  
    -132034.559688351, 
    -1454441.58104013,
  
    -87705.8803012723, 
    -1173951.87151324,
  
    169916.201552955, 
    -2772448.85459782,
  
    -224335.730624953, 
    -1532214.48910552,
  
    -246159.584283012, 
    -1210457.87360091,
  
    291532.63120299, 
    -2367879.88811021,
  
    444985.120484493, 
    -2430186.0451289,
  
    242231.022848571, 
    -1605515.83821897,
  
    11293.9282577625, 
    -1324625.47025355,
  
    -223461.122561186, 
    -1054301.57051493,
  
    -124510.510648811, 
    -1047508.04749632,
  
    -182372.361513255, 
    -2039151.15514534,
  
    254167.529353547, 
    -2484169.93617742,
  
    296954.677827014, 
    -1050311.58389072,
  
    48139.1450644218, 
    -1201051.15269648,
  
    469843.88831142, 
    -2124335.53912032,
  
    269766.876448115, 
    -2466164.45049903,
  
    243244.650476627, 
    -2092150.8476567,
  
    384983.214509501, 
    -1564307.48086196,
  
    -195614.397537858, 
    -1111468.57015512,
  
    457697.055149307, 
    -1791216.76677824,
  
    263451.150888602, 
    -2158083.55208124,
  
    32975.1900275724, 
    -3078660.42218594,
  
    -211536.782757141, 
    -1008988.7000949,
  
    541956.838154933, 
    -2071751.08683451,
  
    118530.217545599, 
    -2598363.0277187,
  
    -160619.607547258, 
    -2670354.42856919,
  
    401404.990048204, 
    -2095936.01392907,
  
    -188378.386715927, 
    -1021420.35637321,
  
    -166219.986914279, 
    -2019788.53017061,
  
    153259.404456401, 
    -2521490.49263858,
  
    -208042.861189015, 
    -1074347.56728906,
  
    205500.894616254, 
    -1582805.46063402,
  
    -4333.02377693533, 
    -1353771.46013622,
  
    391034.881207252, 
    -2236239.81328197,
  
    -108408.831572139, 
    -1457301.80722698,
  
    377769.994050634, 
    -2180093.82266054,
  
    -197182.604171837, 
    -1695923.46737751,
  
    370010.036310497, 
    -2462564.57380652,
  
    -107367.865515646, 
    -1184440.72083149,
  
    46980.7380963933, 
    -1330601.77608204,
  
    -145731.828558434, 
    -1658568.06861993,
  
    -293435.123849041, 
    -1281027.99161158,
  
    302724.653670538, 
    -1845014.56087404,
  
    957.987725184025, 
    -2088103.57236396,
  
    -82213.8692605476, 
    -3140119.32348681,
  
    47161.1645593214, 
    -1176342.49007008,
  
    235550.799460872, 
    -2495332.37442015,
  
    291955.27645244, 
    -2399881.16327738,
  
    -285814.828680165, 
    -1053750.95712609,
  
    -68642.7935884021, 
    -1350161.68551464,
  
    120223.179710297, 
    -2419781.39371525,
  
    -24587.5001732527, 
    -1263222.35146403,
  
    58497.7950173483, 
    -1155771.94197436,
  
    305757.317807243, 
    -1916615.78345423,
  
    158487.370447957, 
    -2350095.77216789,
  
    -264194.975055246, 
    -1178662.1469774,
  
    98819.6711560911, 
    -1981710.89261363,
  
    375711.61106594, 
    -1497944.73880356,
  
    459716.804894248, 
    -1410728.81800095,
  
    485855.211373602, 
    -1760241.128621,
  
    -37055.0931094775, 
    -3070792.6450959,
  
    33232.6648646956, 
    -1352759.43410081,
  
    263586.615019333, 
    -2391617.54896109,
  
    28260.8486396786, 
    -3096107.77561158,
  
    179067.548597284, 
    -2375366.30981703,
  
    -188571.36890161, 
    -1778697.60486185,
  
    -160531.863136307, 
    -2852020.64925544,
  
    83399.1143377826, 
    -2377561.63530107,
  
    400052.772822695, 
    -1510230.66792202,
  
    -249710.313466181, 
    -1058113.60154329,
  
    253293.295431088, 
    -1316175.7067744,
  
    51881.9119296778, 
    -1372464.30662845,
  
    -260600.56698639, 
    -1795825.77386034,
  
    280942.220816244, 
    -1714233.49838976,
  
    -179468.156152233, 
    -1821469.13068435,
  
    231260.757072057, 
    -1564677.26049108,
  
    370165.177372204, 
    -2208619.04746072,
  
    -89193.246849449, 
    -1217019.80907699,
  
    95421.1555174961, 
    -1138046.59847169,
  
    -290210.909889668, 
    -1368023.37975561,
  
    62093.3654112978, 
    -1250640.63595836,
  
    569073.717520117, 
    -1540231.85987997,
  
    279895.336851807, 
    -2337119.13542571,
  
    324933.148367315, 
    -1835382.3730185,
  
    355081.085905086, 
    -2215428.46826378,
  
    -193099.649393767, 
    -2506158.92097258,
  
    446772.200712427, 
    -2099190.8679189,
  
    28579.495404455, 
    -2858173.23437127,
  
    -184218.764067071, 
    -1807355.03813,
  
    465388.41586181, 
    -1803890.09635503,
  
    385757.461930368, 
    -1541472.83723836,
  
    -22895.6621507161, 
    -1325974.21222432,
  
    -49955.722812798, 
    -2859983.56516151,
  
    -169062.392572652, 
    -2381799.56395855,
  
    -198937.0931731, 
    -1800861.85666324,
  
    -14661.6461850226, 
    -1027131.2912839,
  
    351970.777358876, 
    -1535650.88840264,
  
    384912.913245075, 
    -2057652.77107929,
  
    112706.270299012, 
    -1330452.26310989,
  
    84156.6440479159, 
    -1078571.56571105,
  
    -160594.151704685, 
    -2248312.55400777,
  
    -92773.6061254299, 
    -2007851.91280541,
  
    477259.544834189, 
    -1566804.46777282,
  
    201992.156234427, 
    -1553914.80799103,
  
    3550.10240544039, 
    -1308765.3917671,
  
    125359.815640304, 
    -2091369.56482671,
  
    -57261.4720545133, 
    -1259332.11339636,
  
    39590.5985999595, 
    -1123515.9009271,
  
    353771.497603437, 
    -2106419.19709869,
  
    -149423.661652798, 
    -1423794.01943441,
  
    115419.998289885, 
    -1222808.00670836,
  
    361897.862707436, 
    -2149707.21465124,
  
    -211774.214652724, 
    -1739315.72806829,
  
    -15390.4701471092, 
    -2854925.46918303,
  
    -56549.7170840447, 
    -1785487.51604029,
  
    184953.294173791, 
    -2631208.4491777,
  
    -171852.552713775, 
    -2888176.79842235,
  
    -367655.413944817, 
    -1355407.32799382,
  
    171521.098209591, 
    -2812709.18190619,
  
    43262.2609717935, 
    -2364902.91095739,
  
    -278556.779213375, 
    -1598109.05390879,
  
    56105.0379460175, 
    -1294764.53089928,
  
    -81757.9282750292, 
    -2398855.69068928,
  
    110590.528908799, 
    -2686784.5511866,
  
    227028.294112076, 
    -1926725.57544933,
  
    273225.865305442, 
    -2354354.8814922,
  
    108022.688239518, 
    -2112186.39797911,
  
    -156517.258727011, 
    -1118532.24632644,
  
    -245751.990057465, 
    -1151274.75912418,
  
    -69396.0996054531, 
    -1418687.29703354,
  
    -119132.975066829, 
    -1372856.46858484,
  
    175099.977117867, 
    -2713326.56241875,
  
    41621.3814231419, 
    -2312033.74998453,
  
    407243.366113896, 
    -2231725.88257397,
  
    137090.957557004, 
    -1144656.52319521,
  
    59635.7424356703, 
    -1273370.33945888,
  
    -74508.2039407417, 
    -1228959.50523354,
  
    -227058.987294349, 
    -1670461.97428945,
  
    378901.436317771, 
    -2360730.17256556,
  
    389347.188354399, 
    -2074631.43598181,
  
    17410.5351287348, 
    -1163804.62319747,
  
    321641.594479191, 
    -2421236.75026759,
  
    -96726.8748051699, 
    -1468323.73974271,
  
    -184299.517629117, 
    -2159962.98120676,
  
    -128996.269183527, 
    -1173723.40055705,
  
    -141355.641931218, 
    -2916017.57076221,
  
    -137887.961883451, 
    -1341764.36246895,
  
    335710.648866359, 
    -1964586.63715894,
  
    351512.710177393, 
    -2123685.00582727,
  
    229539.279826378, 
    -2214402.71276186,
  
    -197581.41333727, 
    -1842369.49429609,
  
    371094.476788777, 
    -1161200.21551445,
  
    -90042.6580272268, 
    -1750486.68609905,
  
    208483.583461682, 
    -2611868.86065221,
  
    -147060.185166889, 
    -1459801.74703391,
  
    150726.624725493, 
    -2792950.02156658,
  
    -93675.4569681327, 
    -1189068.70774646,
  
    269226.791182248, 
    -2375290.93501582,
  
    458545.328982192, 
    -2430844.49693156,
  
    -233120.378195378, 
    -1064154.02598145,
  
    -54581.9447129313, 
    -1300270.67405077,
  
    127355.650670133, 
    -2074728.36452712,
  
    44350.2574016354, 
    -1401190.25269068,
  
    -140004.738056471, 
    -3010818.98460738,
  
    325045.623306526, 
    -2478371.03004764,
  
    285702.076777369, 
    -1035644.64799243,
  
    36125.2442093186, 
    -1189274.60030435,
  
    263448.419971232, 
    -2451834.97005267,
  
    37009.62010165, 
    -2380485.21683549,
  
    400473.949089309, 
    -1576381.54728283,
  
    272771.830076017, 
    -1080713.51903728,
  
    468074.905177344, 
    -1781286.36142323,
  
    12423.9757656156, 
    -1022046.37873089,
  
    -175049.512580877, 
    -2678646.15240682,
  
    417539.077259274, 
    -2091474.81468459,
  
    -216511.891210187, 
    -2703793.47903624,
  
    -78154.1452217413, 
    -3117800.44365041,
  
    -178724.404816316, 
    -1489552.6349877,
  
    -290105.749881823, 
    -1475433.5219551,
  
    -190662.37620767, 
    -2832951.92060989,
  
    93640.3823603722, 
    -1113243.40462987,
  
    -299998.714077503, 
    -1397005.17704801,
  
    51023.8077071677, 
    -2432305.78883659,
  
    347721.442507151, 
    -1584653.96247938,
  
    -114531.357361067, 
    -1202580.92578436,
  
    30088.5046172605, 
    -1337376.83192649,
  
    -150825.245717378, 
    -1644387.63810128,
  
    63357.5378142827, 
    -1747205.90236138,
  
    121822.742483847, 
    -1585144.53792034,
  
    -48006.021453824, 
    -2735024.07639821,
  
    -63555.3236971478, 
    -1457029.36606999,
  
    61382.2497690024, 
    -1185532.61839973,
  
    307965.147959844, 
    -2397321.6299541,
  
    224677.468880442, 
    -2631456.54627914,
  
    229868.72216474, 
    -2591606.98972139,
  
    514920.534943227, 
    -1932412.45699148,
  
    -28815.9050992973, 
    -2781272.95272826,
  
    -7893.66266204912, 
    -1263574.09268662,
  
    126077.48175422, 
    -2404797.05493669,
  
    214932.52722824, 
    -2172873.63614427,
  
    -400822.625895047, 
    -1121433.85114601,
  
    -16879.3190653113, 
    -1746118.55935286,
  
    -35264.8551075445, 
    -1468580.40165211,
  
    -124643.142990516, 
    -3003759.04169962,
  
    -138586.266781872, 
    -1436017.75546912,
  
    358644.720348683, 
    -2180223.67975637,
  
    466191.710238512, 
    -1825587.57061735,
  
    -159761.08349047, 
    -2740548.36120016,
  
    -204018.205981658, 
    -1372573.04354864,
  
    -36289.8833551283, 
    -1619700.9318212,
  
    416868.923226407, 
    -1499130.82670569,
  
    -159203.271537309, 
    -2215352.56209474,
  
    -141593.324116017, 
    -1524152.59400877,
  
    230697.042408959, 
    -1310487.03496368,
  
    139843.179714918, 
    -2859491.08679711,
  
    87263.3632274778, 
    -2627139.64584784,
  
    -167323.653173065, 
    -1692975.9007161,
  
    356762.388761258, 
    -2199218.85503422,
  
    107206.299901145, 
    -1148955.45586458,
  
    404275.819545282, 
    -1810619.5014861,
  
    79144.0554625487, 
    -1249398.99678569,
  
    -363259.219648233, 
    -1461325.52176117,
  
    -107904.347463196, 
    -2673129.15478504,
  
    260018.307347385, 
    -1879656.40565983,
  
    350446.538244261, 
    -1625072.20189525,
  
    66389.584289699, 
    -1772264.8216832,
  
    305931.99030665, 
    -1068709.76375071,
  
    -179599.038288556, 
    -2973128.53733956,
  
    133580.130062581, 
    -1161787.57002824,
  
    47888.1257116253, 
    -2449843.70607518,
  
    479251.604585636, 
    -1790747.96646017,
  
    97083.0798007573, 
    -2710683.74986074,
  
    -313447.154675126, 
    -1605178.3261813,
  
    -191259.545046386, 
    -1740688.88805916,
  
    -212227.385123593, 
    -1811023.07609872,
  
    123488.291858845, 
    -2539834.25665995,
  
    7272.9845661357, 
    -970428.138720299,
  
    260800.787909039, 
    -2192654.79848367,
  
    40345.5949234557, 
    -1084045.05853702,
  
    -222055.904282248, 
    -1767041.92714597,
  
    221288.068123618, 
    -2415719.0129062,
  
    -168266.168101821, 
    -1724851.16347816,
  
    244718.39483489, 
    -1624646.2826258,
  
    -94352.345781398, 
    -1342853.82257272,
  
    -55857.5531759746, 
    -2787399.0510003,
  
    -309557.261091832, 
    -1326335.03381722,
  
    104699.958409909, 
    -1162845.75558818,
  
    66932.2241921843, 
    -2473833.72420332,
  
    409241.266087628, 
    -2060983.27456036,
  
    -58109.9894780598, 
    -1494614.71967484,
  
    348514.074241251, 
    -2140123.82608489,
  
    -3288.95178220907, 
    -1897545.20827722,
  
    161085.435507945, 
    -2269407.90647356,
  
    -39857.830555191, 
    -1601844.42897566,
  
    -225100.6809214, 
    -1824335.88549759,
  
    -343548.451662017, 
    -1186903.06393152,
  
    -151814.501362441, 
    -2884165.39174597,
  
    19411.7659684552, 
    -1518020.81883901,
  
    -1685.40388907855, 
    -3089932.04493725,
  
    -188155.324452179, 
    -2652640.69773731,
  
    39952.6099357114, 
    -1300688.0805951,
  
    -245630.74307829, 
    -1910213.39049197,
  
    111097.273164438, 
    -1240107.29358136,
  
    -210854.799030644, 
    -1444366.60711208,
  
    -260199.424943524, 
    -1151174.15922403,
  
    -213043.461512157, 
    -2909845.88349818,
  
    281852.762422693, 
    -1690542.27297859,
  
    179660.50986933, 
    -2700203.56633397,
  
    -29525.9933188428, 
    -3056864.906749,
  
    -208411.946798275, 
    -1714069.37576346,
  
    -66080.8798326054, 
    -1212531.56197941,
  
    422274.359819655, 
    -1304819.59142108,
  
    453370.049507853, 
    -2267076.28945735,
  
    405660.053093643, 
    -2072958.0015577,
  
    -100032.064628024, 
    -3018834.66872448,
  
    327861.009435971, 
    -2435746.6202411,
  
    348477.853343095, 
    -1516710.10525593,
  
    499902.025841102, 
    -1697994.38944795,
  
    -155722.902567515, 
    -2361130.16866694,
  
    -253429.500590098, 
    -1583024.49896423,
  
    -75268.2980227616, 
    -1870410.23491718,
  
    294750.714105487, 
    -2185472.36883577,
  
    521723.304974704, 
    -1529014.48462453,
  
    -332793.927745077, 
    -1152699.90890533,
  
    423494.836293606, 
    -2443730.4576161,
  
    130441.76773881, 
    -2454038.49196616,
  
    -113173.43735671, 
    -1766121.18790092,
  
    209664.553135395, 
    -2627613.15006016,
  
    220584.284905885, 
    -1891412.19464274,
  
    132270.279498263, 
    -2797590.63757638,
  
    -99645.031179971, 
    -1204185.54372164,
  
    164792.871926317, 
    -2120270.10923847,
  
    384975.634419029, 
    -1274883.65374691,
  
    21050.6514599944, 
    -1989860.66417495,
  
    -38265.1315616881, 
    -1296427.76903533,
  
    -296260.135267, 
    -1557117.74137763,
  
    27047.0266024822, 
    -1399993.25438059,
  
    -128264.021579468, 
    -3022401.34815127,
  
    331147.51443851, 
    -2465018.63047426,
  
    -139434.619267931, 
    -3160666.57079252,
  
    293596.17338464, 
    -1022053.29389459,
  
    24111.3433542213, 
    -1177498.04791222,
  
    463831.285009056, 
    -2156136.6262169,
  
    256946.581527009, 
    -2437089.60142814,
  
    416225.646199854, 
    -1588659.01509082,
  
    289445.831310248, 
    -1086279.38520503,
  
    25258.649978251, 
    -2106709.28837179,
  
    -135372.048769773, 
    -1729427.64556546,
  
    -132747.295158215, 
    -2655633.45347126,
  
    -218572.891921476, 
    -1548770.82721677,
  
    433673.164470343, 
    -2087013.61544011,
  
    216020.283084302, 
    -2566353.1260944,
  
    282407.871051386, 
    -1507970.49082724,
  
    -184991.173525467, 
    -2022857.51254552,
  
    -273247.47560551, 
    -1624937.42714448,
  
    434921.705778264, 
    -2402024.00624812,
  
    -265653.642257083, 
    -1455760.2050026,
  
    426838.464598721, 
    -1781643.13237201,
  
    -176739.274801237, 
    -2859109.02102808,
  
    378490.612975305, 
    -2234698.52648024,
  
    -121259.874798829, 
    -1484462.92331773,
  
    -44067.1970788064, 
    -3034378.41629203,
  
    78019.5514660794, 
    -2394288.02509278,
  
    -81054.1081587511, 
    -2665584.52997981,
  
    400508.6936284, 
    -1640400.21627821,
  
    -108652.053250428, 
    -1386163.94813386,
  
    -189511.271608938, 
    -3005543.28866167,
  
    95515.1542749351, 
    -1492540.96082928,
  
    235725.080870488, 
    -1108351.68458768,
  
    -190303.281335401, 
    -2894889.83553915,
  
    -226008.796368789, 
    -1897775.66035806,
  
    261233.27660813, 
    -2407917.14430152,
  
    250966.173330907, 
    -2462550.90705833,
  
    238509.412238737, 
    -2619555.65089321,
  
    -140800.289196162, 
    -2056529.66270688,
  
    8800.17704614682, 
    -1263925.83119616,
  
    229821.481374563, 
    -2171653.95839572,
  
    -131614.773560124, 
    -1363608.26665845,
  
    399072.083873845, 
    -1489572.6484479,
  
    38842.8008929675, 
    -1415974.35461144,
  
    4092.53157630286, 
    -1365186.53326211,
  
    345163.011973127, 
    -2172008.06866367,
  
    129710.969775319, 
    -2762058.75570649,
  
    -79509.0716372438, 
    -1815138.35449637,
  
    -175673.079519956, 
    -1672225.53929585,
  
    -125642.56033273, 
    -1825718.60619342,
  
    -79860.2619879327, 
    -1629611.51644077,
  
    -30142.7652768012, 
    -3113432.85308088,
  
    450161.326141053, 
    -2035270.20724667,
  
    91930.7153178815, 
    -2948725.51837011,
  
    696975.69145527, 
    -2095316.12601704,
  
    477637.471884664, 
    -1750764.6791387,
  
    -180057.772750301, 
    -1034317.23010567,
  
    126046.580231469, 
    -1187798.69678103,
  
    343359.600150299, 
    -2189818.66260768,
  
    -80051.1940367928, 
    -1161118.05006003,
  
    250647.001104142, 
    -1923692.63910413,
  
    87471.711634568, 
    -1171213.94753761,
  
    -31430.1946220049, 
    -3087972.28222937,
  
    396353.252521645, 
    -2399213.54017795,
  
    152147.869231091, 
    -1353913.78827848,
  
    349562.105483486, 
    -1604703.72505264,
  
    -423853.466209723, 
    -1138264.8396138,
  
    277283.418080319, 
    -2272305.77043855,
  
    -166478.279925476, 
    -2959343.43120251,
  
    669302.488357685, 
    -2126266.10647082,
  
    -286513.515364118, 
    -1589169.07325685,
  
    -253864.372488296, 
    -1402906.76455536,
  
    355243.366870519, 
    -2072318.75485858,
  
    -237919.166202762, 
    -1767857.45488361,
  
    49015.1567854746, 
    -1385264.64486547,
  
    -84129.7999588294, 
    -2983942.5929848,
  
    -211592.01127349, 
    -1833409.82356303,
  
    -103710.360296755, 
    -2552049.08590575,
  
    231738.683132454, 
    -2277169.60441393,
  
    70097.7658436776, 
    -1145000.41773666,
  
    425303.434149156, 
    -1248266.89098883,
  
    551879.9183297, 
    -1541149.92606466,
  
    89898.6408511076, 
    -2488750.80096405,
  
    431779.886575778, 
    -2181380.2391034,
  
    545405.453675113, 
    -1522644.20515919,
  
    174030.514490705, 
    -2392657.78480159,
  
    -190928.571161609, 
    -1551844.40706194,
  
    -359316.974323214, 
    -1211542.91046881,
  
    66673.6812874672, 
    -1304316.16234526,
  
    -37723.1198290276, 
    -2954528.4672551,
  
    225432.660012423, 
    -1906914.72557339,
  
    -189007.370688402, 
    -2669584.35819302,
  
    -211561.247614337, 
    -2755273.7428373,
  
    82360.2471109197, 
    -3108167.4976059,
  
    -93676.1492282408, 
    -1995927.629486,
  
    421596.681539912, 
    -2255692.39223944,
  
    268572.936519488, 
    -1942809.21814318,
  
    413816.457388754, 
    -1462616.65104202,
  
    467358.36442956, 
    -2364025.4055837,
  
    56889.6350237069, 
    -1083414.70401353,
  
    -57653.5557244748, 
    -1196103.61872529,
  
    368038.217087252, 
    -1695575.67467708,
  
    43062.4774342963, 
    -1152726.41230384,
  
    421972.91757485, 
    -2071284.56467855,
  
    96121.836244399, 
    -1604398.04516863,
  
    318769.565377524, 
    -2447561.97798026,
  
    -124642.02450887, 
    -1188882.84059156,
  
    -91922.8114102642, 
    -2415136.03652506,
  
    -19050.2320692128, 
    -3028328.1112879,
  
    260794.852460852, 
    -2209656.47712461,
  
    402722.923028976, 
    -2357625.59273744,
  
    423525.542100094, 
    -2472068.21259755,
  
    2711.45702655408, 
    -1054926.42389407,
  
    117096.703292449, 
    -2437757.26377737,
  
    -371696.102774852, 
    -1115246.71900378,
  
    149287.225298644, 
    -1982351.07270888,
  
    371668.255298968, 
    -2040144.65378177,
  
    196213.861166382, 
    -1888274.53021558,
  
    -175610.041825715, 
    -1582017.48790758,
  
    264514.132373797, 
    -2132103.56727564,
  
    84751.4194359379, 
    -2779284.13593671,
  
    -231354.371487701, 
    -1157128.0413486,
  
    -403283.726047548, 
    -1404699.65519353,
  
    -32031.2405440521, 
    -1804202.56028305,
  
    -21948.3184104475, 
    -1292584.8640199,
  
    49232.1653121153, 
    -2346532.49288301,
  
    337249.403373506, 
    -2451666.23361389,
  
    282347.764871363, 
    -2319767.65657802,
  
    312424.160587435, 
    -1023110.97075098,
  
    250436.120372095, 
    -2422324.68123919,
  
    -131015.514469788, 
    -2739261.23397362,
  
    238602.064470897, 
    -1742805.39652439,
  
    113187.387647199, 
    -899318.770081004,
  
    47084.5176778141, 
    -2786927.65394086,
  
    -34658.5339836767, 
    -1028474.93197899,
  
    29767.9284370563, 
    -1023332.14769097,
  
    223829.350669195, 
    -2129502.96670023,
  
    4536.13289988753, 
    -2341282.99020299,
  
    498151.010914966, 
    -2054643.38720895,
  
    4454.21801595445, 
    -2531672.13007686,
  
    -61381.3764460226, 
    -2068204.4783434,
  
    95790.9307105364, 
    -1355865.52632177,
  
    129864.220414993, 
    -2377834.23203498,
  
    -140434.750436438, 
    -1931006.34187409,
  
    -168308.038988361, 
    -2043869.44163538,
  
    -184653.481701677, 
    -2913148.9644042,
  
    89824.4179913905, 
    -1203912.87777211,
  
    -205668.733457883, 
    -1912348.2737776,
  
    -28540.8884657744, 
    -2765764.3196904,
  
    25494.0145573509, 
    -1264277.57241876,
  
    279665.403083703, 
    -1305342.46941927,
  
    -188461.842274873, 
    -1385039.14754831,
  
    277071.473939068, 
    -2588677.26572704,
  
    -310324.104415597, 
    -1496990.56075728,
  
    -280893.302656986, 
    -1339579.16333674,
  
    -167237.210855977, 
    -1478912.76485552,
  
    60687.686100418, 
    -1338049.32041756,
  
    49802.1562052021, 
    -2120862.37190994,
  
    346542.604198309, 
    -2158707.25922134,
  
    -102564.681841511, 
    -1402326.79152063,
  
    104857.073576245, 
    -2759728.16902477,
  
    265912.786413347, 
    -2105646.86459798,
  
    -143351.363379984, 
    -2975521.88190711,
  
    -100709.329527657, 
    -1618399.62289298,
  
    -295225.281745393, 
    -1332957.09980449,
  
    -88573.8599682381, 
    -1413925.97239437,
  
    303713.682577305, 
    -1007644.49860851,
  
    558225.118360745, 
    -2118669.12124151,
  
    -9723.17408235443, 
    -1139581.97403848,
  
    187473.770626872, 
    -1326899.88183477,
  
    560465.188228325, 
    -1503292.07185983,
  
    -3766.40426463998, 
    -1984244.83065973,
  
    123256.481582727, 
    -2582948.05584153,
  
    -230048.204968339, 
    -1468338.25395589,
  
    -74870.040258049, 
    -3070074.28676237,
  
    100098.650126158, 
    -1182902.00763608,
  
    405624.568235657, 
    -1350931.44726174,
  
    156951.47647055, 
    -1337623.79034475,
  
    471412.671987683, 
    -2194415.15577216,
  
    435295.612950823, 
    -2213848.7292942,
  
    -77187.8039989129, 
    -960149.770218854,
  
    83107.1220380813, 
    -2796996.12276194,
  
    100866.048577398, 
    -2254759.44859328,
  
    480394.318150249, 
    -1807196.40327633,
  
    239299.63090787, 
    -2481591.39535257,
  
    -220538.719026661, 
    -1725432.64096439,
  
    -253430.827443189, 
    -1771330.32794127,
  
    -230171.105976856, 
    -1866436.56891813,
  
    360279.542032371, 
    -2057687.10630833,
  
    441755.61277412, 
    -2372996.84801774,
  
    -166112.329535759, 
    -1741129.49838875,
  
    453446.638993438, 
    -1775164.00604094,
  
    304475.053765088, 
    -1990648.77132511,
  
    577975.27698828, 
    -2039100.68125376,
  
    -64632.7058166053, 
    -1154824.82446922,
  
    106774.548297021, 
    -1257406.58290938,
  
    213710.771756738, 
    -2276733.76846603,
  
    85351.3504350273, 
    -1155742.6735574,
  
    356308.183868225, 
    -1734674.35410467,
  
    -300383.039547886, 
    -1463855.25025528,
  
    351860.318932786, 
    -2341687.16224491,
  
    -243993.986000595, 
    -1690189.97739865,
  
    434742.969794326, 
    -2165136.31310112,
  
    71580.6666578324, 
    -2835354.90839824,
  
    -369495.43990712, 
    -1199332.81440708,
  
    -106552.92740554, 
    -2655713.58243218,
  
    472513.961725071, 
    -2277024.46104906,
  
    381893.338241876, 
    -1859399.28847154,
  
    -262084.966022424, 
    -1085727.38826502,
  
    -95408.1978568231, 
    -3052263.72906395,
  
    5052.41397039379, 
    -3052003.02932913,
  
    -250195.34149688, 
    -1120120.12455152,
  
    75556.4272286922, 
    -2575350.86148338,
  
    125216.322671824, 
    -2922359.42576861,
  
    -107942.083393916, 
    -1992743.23494885,
  
    -257133.502289755, 
    -1238747.88169579,
  
    -12703.8673345645, 
    -994256.849477032,
  
    -195028.765605778, 
    -1712201.80228815,
  
    -49226.2316163494, 
    -1179675.67547117,
  
    272482.579347446, 
    -1836075.78043778,
  
    30865.8707047279, 
    -1140651.09271708,
  
    -138152.596404659, 
    -2007447.54491021,
  
    309678.121319085, 
    -2459377.33571939,
  
    415433.01463308, 
    -2188040.77408441,
  
    -240950.783953624, 
    -1035662.29170475,
  
    172291.591900014, 
    -1969430.03518294,
  
    -277198.343865524, 
    -1200125.52681073,
  
    -66940.2850811274, 
    -2234552.32688115,
  
    351333.976056836, 
    -1841945.31802281,
  
    20883.810320169, 
    -1052521.14021037,
  
    337937.342445622, 
    -1040260.72181806,
  
    -217430.847798968, 
    -1500737.58077682,
  
    -169398.030005237, 
    -2144332.26203001,
  
    329569.983580036, 
    -1851259.13330195,
  
    -122414.099871036, 
    -1294088.95486616,
  
    -215021.044460939, 
    -1950428.15759261,
  
    -131297.44908038, 
    -2232403.65230367,
  
    305745.376767521, 
    -2127764.15333915,
  
    -5631.50771423514, 
    -1288741.95926251,
  
    133587.488370588, 
    -2776037.37154387,
  
    337961.421967527, 
    -1154294.49131289,
  
    292233.270005294, 
    -2227619.16885112,
  
    238936.894158983, 
    -1759531.5113024,
  
    -120885.153202298, 
    -1802354.2346149,
  
    -133353.094768373, 
    -1746243.97958955,
  
    304819.058460856, 
    -1538016.2594054,
  
    -210484.202776329, 
    -1106127.46714857,
  
    -139146.333057371, 
    -2168556.77930554,
  
    376409.569371702, 
    -2488294.43660966,
  
    131934.276070579, 
    -2359536.03094311,
  
    352683.014395147, 
    -1142565.71689968,
  
    18070.5011841822, 
    -2520038.95632346,
  
    431103.806346408, 
    -1797752.24524455,
  
    -167191.138272758, 
    -1142211.45005116,
  
    357649.946375713, 
    -1173060.69994723,
  
    -72764.9225366169, 
    -3025342.24126392,
  
    -136339.820421505, 
    -3053820.10570149,
  
    456417.891036039, 
    -2136243.26929372,
  
    -260392.952697743, 
    -1202156.42584157,
  
    -431604.509902741, 
    -1314525.98975835,
  
    -72579.8351159461, 
    -1191792.92738907,
  
    -133660.066820528, 
    -3036882.69375381,
  
    -169402.986554564, 
    -2912678.9689119,
  
    84180.8471136991, 
    -1236380.80496284,
  
    271966.491458689, 
    -2484108.92752824,
  
    -188929.263382599, 
    -1907956.40982997,
  
    -262968.143096624, 
    -1388448.82464395,
  
    -108422.632700421, 
    -2057331.40170608,
  
    42187.851810522, 
    -1264629.31118634,
  
    -44591.5908350703, 
    -2585840.88089345,
  
    -161013.168758132, 
    -1373255.66721542,
  
    269190.925542158, 
    -951212.43151803,
  
    7483.67772606654, 
    -2602287.07610393,
  
    -7472.60478577426, 
    -1969690.81621875,
  
    -210947.737002195, 
    -1994555.73888201,
  
    -225155.797062637, 
    -1808288.50060662,
  
    -43405.3014378617, 
    -2943003.07593019,
  
    -488.19024537437, 
    -3113856.49031568,
  
    90354.7529378385, 
    -2965926.25612081,
  
    477632.327426707, 
    -1845377.75680896,
  
    -85789.5532653301, 
    -1479229.8228246,
  
    432999.518677607, 
    -2420586.75108892,
  
    576133.019611719, 
    -1512470.15641593,
  
    -191032.545123172, 
    -2867118.39163338,
  
    539.014781406914, 
    -2105537.34472802,
  
    -30197.6331347369, 
    -1942243.74860027,
  
    60181.611359625, 
    -2815618.81090201,
  
    142560.376099123, 
    -1102255.73585701,
  
    494828.864754878, 
    -1802278.49043303,
  
    -241715.459869599, 
    -1747050.09024577,
  
    149933.860828745, 
    -936114.34579198,
  
    272677.361139816, 
    -1064818.40228561,
  
    16093.8045267766, 
    -1385153.66057025,
  
    49362.1857862104, 
    -2104752.28629073,
  
    -86399.2378976354, 
    -2691462.40352427,
  
    134857.273944503, 
    -2810946.69081575,
  
    411066.295757881, 
    -1542223.79380918,
  
    -70772.8409457939, 
    -1170373.57184867,
  
    71224.2838324307, 
    -1119701.45835878,
  
    102458.932069953, 
    -1274680.15221776,
  
    72049.0873340201, 
    -2869237.59983423,
  
    -176587.157528148, 
    -1645452.68952607,
  
    -274859.032023768, 
    -1442007.32108924,
  
    410730.520860246, 
    -2464529.75788693,
  
    437706.055725928, 
    -2148892.38929577,
  
    379950.647386432, 
    -2250783.992463,
  
    30615.5475554687, 
    -2840314.14439766,
  
    23053.96053334, 
    -1750046.97075159,
  
    434552.410387411, 
    -1509191.1053722,
  
    30845.9438089876, 
    -1312979.38131485,
  
    69634.150321348, 
    -2852718.79208173,
  
    -62636.5353901341, 
    -2769490.4339654,
  
    -193304.418041778, 
    -2730838.95604384,
  
    -246755.870010558, 
    -1089948.75484353,
  
    280385.424534519, 
    -2065502.67762789,
  
    -12000.9401467111, 
    -3074988.32949666,
  
    354192.18436443, 
    -1359506.55668148,
  
    67715.2257987948, 
    -1075948.40899648,
  
    -40798.9075082297, 
    -1163247.73221706,
  
    277778.28272799, 
    -1851702.32754618,
  
    18669.2664301917, 
    -1128575.7728723,
  
    354043.102835497, 
    -2244427.27500185,
  
    72550.2611951717, 
    -1208354.99481906,
  
    300586.677260652, 
    -2471192.69345848,
  
    402049.226166951, 
    -2178457.38551819,
  
    -177748.295136262, 
    -2777002.27074957,
  
    162528.219578257, 
    -2620452.3387008,
  
    -138541.619133011, 
    -993214.544400501,
  
    54975.7052395826, 
    -1869154.53754808,
  
    154884.781285695, 
    -1886645.61094942,
  
    191464.280772064, 
    -1008978.67854555,
  
    366102.337181609, 
    -2028338.63084122,
  
    122120.078834325, 
    -1205015.83520276,
  
    -134439.500925597, 
    -2250912.82020163,
  
    363273.703000878, 
    -1748876.96391593,
  
    10685.3054370008, 
    -1284899.05424708,
  
    -53754.5256546383, 
    -1166579.32068057,
  
    349826.948563987, 
    -1978677.90447123,
  
    474836.50560659, 
    -2092208.43054717,
  
    118007.124499446, 
    -987145.697065475,
  
    -75329.8447430995, 
    -1444946.00969775,
  
    -439356.788194462, 
    -1271982.32717442,
  
    -31608.939054731, 
    -996164.57780223,
  
    -208254.588563992, 
    -1591266.90205571,
  
    148115.735233021, 
    -2495855.51626931,
  
    459493.428280567, 
    -1923240.0953751,
  
    -284069.113095863, 
    -1419054.00452954,
  
    401691.390042364, 
    -1790885.30685593,
  
    -66665.712009243, 
    -2300775.63471118,
  
    -141315.934374039, 
    -1470598.47146601,
  
    131817.766692888, 
    -2873951.57295756,
  
    -198423.317853421, 
    -2033455.10718396,
  
    -150562.785104924, 
    -3040012.56414955,
  
    72166.9462585784, 
    -1224604.2525707,
  
    313156.12141591, 
    -2408989.29482956,
  
    137908.012805652, 
    -2313353.6372601,
  
    597133.556506003, 
    -2159361.54101286,
  
    -173755.703502156, 
    -2644987.08488107,
  
    -197717.472580733, 
    -1479078.59997196,
  
    -110454.809429712, 
    -2892098.02065715,
  
    460966.181463077, 
    -1318241.90968721,
  
    -238355.620366795, 
    -1815225.7702117,
  
    13716.6484662527, 
    -916555.675197524,
  
    -113159.991558612, 
    -1169632.10679717,
  
    -28540.3615900481, 
    -2942124.67803325,
  
    379932.077387129, 
    -1191095.96638138,
  
    -199413.007533279, 
    -1457074.67529627,
  
    298309.865881564, 
    -2168002.85098835,
  
    282956.866832911, 
    -2385434.68985026,
  
    -308856.35445768, 
    -1583088.08440186,
  
    27682.1305475161, 
    -2760813.43609689,
  
    -110467.084233997, 
    -1715353.00061495,
  
    -224903.12385411, 
    -1751436.40421684,
  
    431853.203671975, 
    -1537218.98349324,
  
    -137752.538271456, 
    -2807953.51942687,
  
    19923.1427400391, 
    -2773367.46149237,
  
    -303081.014395739, 
    -1131283.90681529,
  
    567456.29865403, 
    -2232793.54769493,
  
    440702.100971436, 
    -2132467.76865227,
  
    -258475.06695951, 
    -1876686.94771,
  
    418287.42838674, 
    -1519951.68257491,
  
    -145649.29212085, 
    -1307825.89391538,
  
    370390.200410916, 
    -1485158.0709699,
  
    -98931.4535997581, 
    -1977795.32203217,
  
    -135517.696355456, 
    -1990932.28216887,
  
    554194.346218936, 
    -2047039.77342521,
  
    -168832.436214495, 
    -1423970.47035346,
  
    -81786.1124425425, 
    -2944280.63604516,
  
    -32371.5834001157, 
    -1146819.78896296,
  
    86335.1928408139, 
    -1219492.58895198,
  
    291495.233202226, 
    -2483008.05119753,
  
    388665.437442774, 
    -2168873.99449691,
  
    -57212.6100194664, 
    -1769276.65145021,
  
    136707.454329702, 
    -1843456.0921776,
  
    -18911.1587137596, 
    -3009912.9705982,
  
    656062.03512223, 
    -2217229.2335624,
  
    -2958.27143450601, 
    -2244772.19677985,
  
    357012.703675528, 
    -2426326.25992036,
  
    27002.1185882344, 
    -1281056.14923166,
  
    -47486.4696439081, 
    -1150706.64158919,
  
    291019.876706738, 
    -2415847.72825393,
  
    402130.302328509, 
    -1613658.12187171,
  
    -152312.607782066, 
    -1809652.31791012,
  
    -411314.735977162, 
    -1309965.25694156,
  
    116948.285674441, 
    -1313822.41743523,
  
    -141560.835813337, 
    -1564607.60153523,
  
    283456.202029572, 
    -1289033.99551586,
  
    -517669.853120274, 
    -1208333.44049211,
  
    -181370.907178542, 
    -2990614.47983827,
  
    60153.0456614973, 
    -1212827.70263359,
  
    461202.78731995, 
    -2114629.57269424,
  
    224262.701528291, 
    -2112253.50653861,
  
    312816.14905608, 
    -2474781.86188208,
  
    25195.2151986743, 
    -1219135.09586513,
  
    14265.1883850089, 
    -1248995.58871286,
  
    910.117445646081, 
    -1248714.196329,
  
    303458.706878373, 
    -2444867.47065601,
  
    278858.32076457, 
    -2454349.09521496,
  
    272638.905807761, 
    -2439839.22524148,
  
    36297.5986486253, 
    -2396813.6271965,
  
    381156.419609304, 
    -1584475.7619147,
  
    401302.125708912, 
    -1595019.83457728,
  
    528624.778515938, 
    -1931705.91205638,
  
    -27560.7091470259, 
    -2794582.80778312,
  
    11309.3403785698, 
    -1211928.46985322,
  
    -27797.6206626182, 
    -1236585.90516931,
  
    -47701.5789212004, 
    -1209597.71519699,
  
    127970.849857093, 
    -2391315.64361488,
  
    -120284.789113107, 
    -1439869.50116235,
  
    289304.674495717, 
    -1066764.08314717,
  
    97605.4337601426, 
    -2698358.6198612,
  
    -229410.255079364, 
    -1794811.48553766,
  
    -223089.201875714, 
    -1780790.78496621,
  
    -51794.2918506582, 
    -1505934.51319669,
  
    123007.919718597, 
    -2788035.15285207,
  
    7758.36286611733, 
    -1181219.16512407,
  
    -24947.5964291731, 
    -1188661.39192467,
  
    -24571.3458266078, 
    -1166810.31311113,
  
    -12557.4476845845, 
    -1178586.86330625,
  
    450768.670754547, 
    -2152514.51143888,
  
    273983.228018372, 
    -2426468.66619758,
  
    421434.830559239, 
    -1571512.33970035,
  
    277948.244485576, 
    -1096873.2737713,
  
    419418.120776915, 
    -1767015.16250628,
  
    -163619.455313052, 
    -1679347.66808968,
  
    -169808.14016984, 
    -1042511.19523155,
  
    447783.977576907, 
    -2168586.74505116,
  
    68144.0119464864, 
    -1091014.55012471,
  
    260834.525553013, 
    -2222785.02188412,
  
    -175751.086928943, 
    -2055034.5122407,
  
    -174165.198662327, 
    -1467370.86859514,
  
    64992.9291515771, 
    -1353151.16952448,
  
    105153.17409594, 
    -2746273.23936003,
  
    4473.04630293694, 
    -1134078.8746829,
  
    573090.464525216, 
    -1498144.38159072,
  
    -255979.310436627, 
    -1756997.05197898,
  
    418396.095912663, 
    -2171796.85325023,
  
    168215.579469233, 
    -1956964.39257167,
  
    6123.32319213978, 
    -2513337.70674617,
  
    12305.7683410976, 
    -3111243.89350417,
  
    504666.785019562, 
    -1810316.76688557,
  
    149693.598304323, 
    -922664.176406716,
  
    -286785.334605733, 
    -1433295.21809827,
  
    405012.309643516, 
    -2162213.46197091,
  
    414683.76823762, 
    -2150670.88415866,
  
    35379.5484866149, 
    -2827874.75447853,
  
    43275.8679836303, 
    -2841704.0944428,
  
    305219.484044921, 
    -2487365.74150776,
  
    386119.536197342, 
    -2117516.41163776,
  
    387816.802401666, 
    -2151754.80365598,
  
    412986.502033326, 
    -2116432.49214047,
  
    3470.18026948382, 
    -1335741.76520054,
  
    329144.616142944, 
    -2384172.03810121,
  
    351724.964751191, 
    -2394658.8160287,
  
    -69203.2488696528, 
    -1432487.35868566,
  
    132401.151921222, 
    -2439558.43785173,
  
    -47931.6421681711, 
    -1281570.64473015,
  
    -57814.3664295476, 
    -1229311.24645611,
  
    225611.735820808, 
    -2159214.67073627,
  
    491005.3668252, 
    -1814155.42171282,
  
    -214971.01550994, 
    -1792572.14407207,
  
    96461.2833787248, 
    -1068087.39815162,
  
    314429.109836925, 
    -1051672.2664268,
  
    -134805.839918593, 
    -1716778.17603114,
  
    451728.751858062, 
    -1515322.34944589,
  
    446746.903330097, 
    -1569883.24547675,
  
    46074.8287408167, 
    -1234938.56881524,
  
    60407.5887686232, 
    -1127925.61292952,
  
    427603.062532382, 
    -2120290.51888662,
  
    430638.113759398, 
    -2103652.06961841,
  
    52598.9509003117, 
    -1048851.52303751,
  
    -190794.462743803, 
    -1753049.87986494,
  
    397743.85312878, 
    -2217919.4721315,
  
    -289644.332413081, 
    -1223301.60786284,
  
    -78109.3340061698, 
    -1275549.34843705,
  
    372749.641152579, 
    -2084687.54829668,
  
    27491.3418192236, 
    -1091276.35606894,
  
    -153322.213431376, 
    -1448540.95020008,
  
    435835.568977706, 
    -1554385.25076517,
  
    460529.921953637, 
    -1577761.12408587,
  
    174949.407148405, 
    -2547147.6480675,
  
    17245.7351549697, 
    -1146659.06605892,
  
    -11182.5680539519, 
    -1156193.93437914,
  
    312550.150420746, 
    -2433052.10800679,
  
    412875.779056391, 
    -1627040.18410362,
  
    374818.56822111, 
    -2134177.71597907,
  
    214306.17350145, 
    -2204131.83848517,
  
    222906.011914868, 
    -2607840.11242526,
  
    -232205.953257406, 
    -1044981.93110984,
  
    -215751.994201111, 
    -1064324.57038754,
  
    -174296.174213769, 
    -2029469.84265799,
  
    304800.73476904, 
    -1036515.54755224,
  
    28469.6588583043, 
    -1232488.49465937,
  
    280631.054825177, 
    -2474586.25084829,
  
    398024.755262708, 
    -1553265.63856308,
  
    263982.639434209, 
    -2145093.56239152,
  
    -199957.584478501, 
    -1015204.53068908,
  
    -13614.3452898366, 
    -1339872.83766582,
  
    373967.583643444, 
    -2194356.43900122,
  
    43466.6741450685, 
    -1315644.92956608,
  
    -34960.8449590816, 
    -1250549.65532038,
  
    -41120.5291763878, 
    -1229662.98522367,
  
    -15109.5036857126, 
    -1275982.15781829,
  
    -242878.181895497, 
    -1802057.138461,
  
    67130.1546074268, 
    -1237622.44439355,
  
    -30580.3980837169, 
    -1311200.99075884,
  
    -1118.83605016511, 
    -1024588.83881895,
  
    -9199.10787348858, 
    -1300675.12912101,
  
    -60201.2778345692, 
    -1243731.93075309,
  
    347090.044900572, 
    -2093035.47076046,
  
    190463.059475782, 
    -2619937.23731524,
  
    -275902.127280427, 
    -1611523.24175415,
  
    -235526.487745969, 
    -1680325.97720058,
  
    470302.834016499, 
    -2423152.21972213,
  
    -47695.7378014511, 
    -1315288.24787996,
  
    30660.2284764853, 
    -1204204.84821375,
  
    9713.89975032844, 
    -1233854.29725832,
  
    297239.291921579, 
    -2430357.60068251,
  
    294268.221299865, 
    -2456863.21792221,
  
    64873.5598244785, 
    -1759735.36215132,
  
    60767.6478442669, 
    -1199180.16174417,
  
    17710.3418663979, 
    -1194713.25888272,
  
    -17845.6416623363, 
    -1250079.99892796,
  
    1395.82138747398, 
    -1274236.57346685,
  
    141205.675469968, 
    -2408764.5030034,
  
    -410726.475178627, 
    -1111130.10436491,
  
    129813.353919513, 
    -1174793.13353365,
  
    -299980.335019622, 
    -1597173.69971908,
  
    -274796.159496763, 
    -1148437.361258,
  
    -171326.067265353, 
    -2364904.48503653,
  
    -41300.5771753186, 
    -1192382.50668151,
  
    243250.594472792, 
    -2438830.15972199,
  
    46425.79886336, 
    -1426247.91937784,
  
    -30786.4809188817, 
    -3100702.57023919,
  
    419452.560606733, 
    -1263187.61440941,
  
    265213.458295078, 
    -2118875.21729336,
  
    -164079.508104303, 
    -1491268.45086664,
  
    -132397.170572977, 
    -2965217.33594126,
  
    -78195.3566691598, 
    -1405548.4679486,
  
    104214.029656655, 
    -2241058.03902152,
  
    -239851.435387105, 
    -1859741.89787564,
  
    400569.534851636, 
    -2191663.95186031,
  
    -144478.89837656, 
    -1740092.98367228,
  
    -73732.5790291914, 
    -3012548.7530128,
  
    422242.575729971, 
    -2410364.69293141,
  
    49155.1804017803, 
    -2091377.08704111,
  
    427692.933506031, 
    -2141569.32776201,
  
    166559.584094967, 
    -2607120.22715106,
  
    386968.169299509, 
    -2134635.6076469,
  
    399128.701207724, 
    -2108414.85278603,
  
    -153783.128049995, 
    -3018537.81966202,
  
    -192194.338930493, 
    -1518968.61043366,
  
    -31614.829016934, 
    -1277727.73971471,
  
    49842.3198780133, 
    -1359505.09576783,
  
    -173625.7418973, 
    -1410888.16371277,
  
    465981.934398974, 
    -1945343.12956045,
  
    -201861.663565168, 
    -1788858.82210037,
  
    322163.849860606, 
    -1038071.95875843,
  
    -182885.164491616, 
    -1840727.83169286,
  
    47106.9870316365, 
    -1217994.86198337,
  
    355778.888063557, 
    -2442482.06160359,
  
    -214910.308863625, 
    -1561508.16626483,
  
    133874.284996653, 
    -2345669.1945546,
  
    -414627.233693185, 
    -1257885.041526,
  
    95089.9890919102, 
    -2801473.52778395,
  
    294252.496049756, 
    -2198084.94869241,
  
    230046.091212045, 
    -2185906.99976088,
  
    391144.789715753, 
    -2387665.30021222,
  
    -126647.217243592, 
    -1469452.25217893,
  
    -174387.468067688, 
    -2661497.56709384,
  
    -166832.68138162, 
    -2007387.16502844,
  
    203746.525554358, 
    -1568360.13554004,
  
    299123.804125773, 
    -1832751.90483149,
  
    227518.739681973, 
    -1550382.55493669,
  
    385663.005203646, 
    -2043288.07566508,
  
    197308.923654593, 
    -2629410.79961894,
  
    -178253.019662759, 
    -2900662.88167133,
  
    400825.967928108, 
    -2142653.24971435,
  
    16779.342443372, 
    -1336559.29856351,
  
    -14761.9686189017, 
    -1228366.76023597,
  
    -26847.6141354754, 
    -1220611.06841146,
  
    -222733.754349616, 
    -1074662.02445759,
  
    341094.350680523, 
    -2402002.7484113,
  
    -6819.12925281876, 
    -1200294.93101796,
  
    -47581.063722835, 
    -1247140.79452228,
  
    416250.55960504, 
    -1556868.06836933,
  
    247108.383061391, 
    -2450690.53720173,
  
    399977.334825954, 
    -2125534.05370525,
  
    288048.804404112, 
    -2442353.35311684,
  
    -63020.4890566502, 
    -1278559.99916764,
  
    -241420.541261277, 
    -1783070.90673947,
  
    377463.432752753, 
    -2159730.14518363,
  
    359919.841928079, 
    -2088861.5108851,
  
    413835.135393511, 
    -2133551.69060462,
  
    -143606.075866638, 
    -3027815.57253516,
  
    461039.534187367, 
    -1558387.68355506,
  
    -1712.1024649029, 
    -1168706.55097911,
  
    -253590.547393356, 
    -1807518.85375945,
  
    29653.9307740314, 
    -1250438.93327848,
  
    -1726.31412016385, 
    -1220147.61504459,
  
    -25897.6051533073, 
    -1204636.23139557,
  
    361666.320003668, 
    -2137150.771161,
  
    57118.5695920168, 
    -1227808.65331747,
  
    376140.999388439, 
    -2146953.9319379,
  
    -66959.623460413, 
    -1291336.78911692,
  
    -13811.9593787037, 
    -1212391.9256751,
  
    -148518.141257892, 
    -927096.472804295,
  
    -145924.552917179, 
    -919442.668323767,
  
    -593007.1400445, 
    -1373157.95499468,
  
    -243026.481598873, 
    -3006510.4402062,
  
    -251605.304691925, 
    -3007926.76397332,
  
    812800.481224708, 
    -2029554.24720719,
  
    551988.065703701, 
    -1803374.50238612,
  
    527480.109611981, 
    -2344326.22809166,
  
    578684.207954812, 
    -1833291.24517149,
  
    591474.340634011, 
    -1836854.61248345,
  
    579500.112490506, 
    -1403270.16496941,
  
    515702.484221326, 
    -1088502.05803231,
  
    511947.073248662, 
    -1079961.30742867,
  
    505315.707631775, 
    -1086016.36917192,
  
    785140.460503185, 
    -2079447.03008274,
  
    633422.06425264, 
    -1581194.31982653,
  
    629534.327187448, 
    -1573358.50423487,
  
    567513.837406947, 
    -1866773.91920444,
  
    489809.039829813, 
    -1151970.97826282,
  
    -249591.560341304, 
    -2892780.31839919,
  
    47820.3591706862, 
    -858841.51051191,
  
    544741.114808772, 
    -1671505.77871744,
  
    531317.560443355, 
    -1671342.36241007,
  
    572129.878205254, 
    -1817716.30286775,
  
    -84748.1976712063, 
    -910344.196727883,
  
    -85023.7775194824, 
    -919730.278581974,
  
    124613.187858324, 
    -3103580.33121491,
  
    130805.030796487, 
    -3107794.78436472,
  
    90149.7106894431, 
    -3177526.51726136,
  
    207237.580853052, 
    -2852767.39219661,
  
    283109.91014316, 
    -2651371.886254,
  
    336702.345346114, 
    -2561219.11216479,
  
    549182.258774561, 
    -1914680.5323359,
  
    526554.881696154, 
    -1740842.30628323,
  
    679319.144686799, 
    -2219338.68210279,
  
    -262041.479192898, 
    -1923973.37021481,
  
    276451.123018265, 
    -932766.292352424,
  
    -246311.05490594, 
    -2651140.42645688,
  
    -235717.050623179, 
    -1972068.491574,
  
    160301.29657002, 
    -879569.753803044,
  
    168723.703738361, 
    -874705.265729038,
  
    593495.077340233, 
    -1868946.7522172,
  
    584729.483664223, 
    -1871183.27044853,
  
    156868.121564966, 
    -886230.472844777,
  
    66077.4897556385, 
    -841594.036383364,
  
    68861.9777791475, 
    -848563.878589684,
  
    10527.7035558456, 
    -3166161.1876335,
  
    582344.175316364, 
    -1620241.27741493,
  
    -83956.6879944971, 
    -927880.529395933,
  
    -80191.2370067825, 
    -939102.548437344,
  
    -156720.72580318, 
    -935926.248296663,
  
    651897.025833008, 
    -1593908.78141827,
  
    641418.427840558, 
    -1588238.05013781,
  
    -479716.323360212, 
    -1407231.07774586,
  
    550824.807809979, 
    -1676989.21293295,
  
    600057.887975449, 
    -2277898.99186964,
  
    512705.099691944, 
    -1357582.89251946,
  
    492489.481718792, 
    -1342656.39330972,
  
    500066.078703513, 
    -1344134.63994944,
  
    -246862.853076102, 
    -1963845.2805743,
  
    540746.864479175, 
    -1304286.32883775,
  
    765740.132688, 
    -2120130.37783302,
  
    -236050.719991169, 
    -3002573.17740333,
  
    -257750.194429692, 
    -3012839.75461722,
  
    -160134.702080425, 
    -3125651.44361157,
  
    557814.000747449, 
    -1674093.61067516,
  
    620887.815662721, 
    -1573305.67108534,
  
    613573.263315598, 
    -1575431.72379944,
  
    -319310.650530788, 
    -1044224.33501309,
  
    -524362.98951776, 
    -1414090.12298943,
  
    -517727.434333712, 
    -1410361.78175851,
  
    -472841.862700287, 
    -1278964.94474706,
  
    593402.124214133, 
    -2271870.11554207,
  
    481883.152256224, 
    -1336745.74442852,
  
    488510.945687472, 
    -1329754.72811001,
  
    551467.714796272, 
    -1330410.29865276,
  
    765220.301369214, 
    -2110095.77567314,
  
    745600.492587742, 
    -2154822.71240745,
  
    570901.539661809, 
    -2077233.4493075,
  
    592797.302546144, 
    -2039058.21595414,
  
    252709.15172009, 
    -911893.078177904,
  
    -218394.601319314, 
    -2941701.60740137,
  
    577184.051742036, 
    -1866195.38928562,
  
    55384.399488186, 
    -859232.62111609,
  
    562294.111234805, 
    -1647092.61682083,
  
    134077.247869996, 
    -3110046.1154575,
  
    211286.189705627, 
    -2804600.06802987,
  
    -268184.86360689, 
    -2902906.20257121,
  
    -546746.43437222, 
    -1395568.83757297,
  
    505749.666344389, 
    -1354483.06578604,
  
    485443.808618241, 
    -1346609.95720863,
  
    550274.554192431, 
    -1321774.04951451,
  
    -237488.763831075, 
    -2651034.38432199,
  
    564994.217509373, 
    -2062655.44867261,
  
    580427.847184576, 
    -1851035.35811893,
  
    531474.373375532, 
    -1766206.42987563,
  
    97526.6052949081, 
    -3020538.2508376,
  
    605880.770937027, 
    -1635043.13366869,
  
    600634.995389901, 
    -1628581.23534773,
  
    -249323.785652818, 
    -1930795.41892682,
  
    495774.699043105, 
    -1291950.41485203,
  
    -218273.935077366, 
    -2776804.85242306,
  
    585099.914806698, 
    -1974145.91409993,
  
    94415.4449319034, 
    -860561.814283983,
  
    1598.00427734903, 
    -894178.053894874,
  
    9053.5754574886, 
    -895395.401488985,
  
    538811.211607869, 
    -1695734.80658933,
  
    -81128.0078016883, 
    -947633.877320175,
  
    591780.661320064, 
    -1626222.91062403,
  
    53563.9210653029, 
    -3239100.86679958,
  
    118198.587627829, 
    -3156798.41991678,
  
    607660.110191382, 
    -1589816.29169027,
  
    600827.180756676, 
    -1585659.1518606,
  
    -268943.667079332, 
    -1016423.27539622,
  
    116134.552603853, 
    -3122873.18164566,
  
    121007.584193571, 
    -3129241.08731521,
  
    495907.65490353, 
    -1324727.61294023,
  
    264833.700010829, 
    -901011.391931257,
  
    259671.241507911, 
    -907438.811458146,
  
    125803.949664276, 
    -3158243.83513511,
  
    -511227.572924795, 
    -1405264.13693297,
  
    795106.49350194, 
    -2034839.28457689,
  
    739771.934942861, 
    -2180398.06278457,
  
    795331.823644945, 
    -2058849.25113685,
  
    789400.795007781, 
    -2065634.0907815,
  
    557627.871660767, 
    -1929637.43844612,
  
    35657.2830666926, 
    -3247189.7673356,
  
    -153702.238552524, 
    -943316.97439178,
  
    202722.098867646, 
    -895201.216008158,
  
    151170.565068844, 
    -2932163.5775673,
  
    -519495.560050131, 
    -1236106.00864367,
  
    802965.320179788, 
    -2033487.54773535,
  
    -235412.768588272, 
    -2360147.87297206,
  
    722264.964597462, 
    -2046358.96120813,
  
    132094.132866408, 
    -876899.073613287,
  
    -181113.318791924, 
    -3086678.7412297,
  
    -85101.4019456898, 
    -902337.722171635,
  
    135713.724672627, 
    -3098304.01047402,
  
    543200.698385186, 
    -1313759.6368711,
  
    -425601.082066204, 
    -1429202.68196879,
  
    -245433.921586739, 
    -2700373.66330056,
  
    -212029.351647646, 
    -2811750.62368031,
  
    38212.2211017756, 
    -3239604.53614449 ;

 grid.cells.index = 
    1, 
    2, 
    3, 
    4, 
    5, 
    6, 
    7, 
    8, 
    9, 
    10, 
    11, 
    12, 
    13, 
    14, 
    15, 
    16, 
    17, 
    18, 
    19, 
    20, 
    21, 
    22, 
    23, 
    24, 
    25, 
    26, 
    27, 
    28, 
    29, 
    30, 
    31, 
    32, 
    33, 
    34, 
    35, 
    36, 
    37, 
    38, 
    39, 
    40, 
    41, 
    42, 
    43, 
    44, 
    45, 
    46, 
    47, 
    48, 
    49, 
    50, 
    51, 
    52, 
    53, 
    54, 
    55, 
    56, 
    57, 
    58, 
    59, 
    60, 
    61, 
    62, 
    63, 
    64, 
    65, 
    66, 
    67, 
    68, 
    69, 
    70, 
    71, 
    72, 
    73, 
    74, 
    75, 
    76, 
    77, 
    78, 
    79, 
    80, 
    81, 
    82, 
    83, 
    84, 
    85, 
    86, 
    87, 
    88, 
    89, 
    90, 
    91, 
    92, 
    93, 
    94, 
    95, 
    96, 
    97, 
    98, 
    99, 
    100, 
    101, 
    102, 
    103, 
    104, 
    105, 
    106, 
    107, 
    108, 
    109, 
    110, 
    111, 
    112, 
    113, 
    114, 
    115, 
    116, 
    117, 
    118, 
    119, 
    120, 
    121, 
    122, 
    123, 
    124, 
    125, 
    126, 
    127, 
    128, 
    129, 
    130, 
    131, 
    132, 
    133, 
    134, 
    135, 
    136, 
    137, 
    138, 
    139, 
    140, 
    141, 
    142, 
    143, 
    144, 
    145, 
    146, 
    147, 
    148, 
    149, 
    150, 
    151, 
    152, 
    153, 
    154, 
    155, 
    156, 
    157, 
    158, 
    159, 
    160, 
    161, 
    162, 
    163, 
    164, 
    165, 
    166, 
    167, 
    168, 
    169, 
    170, 
    171, 
    172, 
    173, 
    174, 
    175, 
    176, 
    177, 
    178, 
    179, 
    180, 
    181, 
    182, 
    183, 
    184, 
    185, 
    186, 
    187, 
    188, 
    189, 
    190, 
    191, 
    192, 
    193, 
    194, 
    195, 
    196, 
    197, 
    198, 
    199, 
    200, 
    201, 
    202, 
    203, 
    204, 
    205, 
    206, 
    207, 
    208, 
    209, 
    210, 
    211, 
    212, 
    213, 
    214, 
    215, 
    216, 
    217, 
    218, 
    219, 
    220, 
    221, 
    222, 
    223, 
    224, 
    225, 
    226, 
    227, 
    228, 
    229, 
    230, 
    231, 
    232, 
    233, 
    234, 
    235, 
    236, 
    237, 
    238, 
    239, 
    240, 
    241, 
    242, 
    243, 
    244, 
    245, 
    246, 
    247, 
    248, 
    249, 
    250, 
    251, 
    252, 
    253, 
    254, 
    255, 
    256, 
    257, 
    258, 
    259, 
    260, 
    261, 
    262, 
    263, 
    264, 
    265, 
    266, 
    267, 
    268, 
    269, 
    270, 
    271, 
    272, 
    273, 
    274, 
    275, 
    276, 
    277, 
    278, 
    279, 
    280, 
    281, 
    282, 
    283, 
    284, 
    285, 
    286, 
    287, 
    288, 
    289, 
    290, 
    291, 
    292, 
    293, 
    294, 
    295, 
    296, 
    297, 
    298, 
    299, 
    300, 
    301, 
    302, 
    303, 
    304, 
    305, 
    306, 
    307, 
    308, 
    309, 
    310, 
    311, 
    312, 
    313, 
    314, 
    315, 
    316, 
    317, 
    318, 
    319, 
    320, 
    321, 
    322, 
    323, 
    324, 
    325, 
    326, 
    327, 
    328, 
    329, 
    330, 
    331, 
    332, 
    333, 
    334, 
    335, 
    336, 
    337, 
    338, 
    339, 
    340, 
    341, 
    342, 
    343, 
    344, 
    345, 
    346, 
    347, 
    348, 
    349, 
    350, 
    351, 
    352, 
    353, 
    354, 
    355, 
    356, 
    357, 
    358, 
    359, 
    360, 
    361, 
    362, 
    363, 
    364, 
    365, 
    366, 
    367, 
    368, 
    369, 
    370, 
    371, 
    372, 
    373, 
    374, 
    375, 
    376, 
    377, 
    378, 
    379, 
    380, 
    381, 
    382, 
    383, 
    384, 
    385, 
    386, 
    387, 
    388, 
    389, 
    390, 
    391, 
    392, 
    393, 
    394, 
    395, 
    396, 
    397, 
    398, 
    399, 
    400, 
    401, 
    402, 
    403, 
    404, 
    405, 
    406, 
    407, 
    408, 
    409, 
    410, 
    411, 
    412, 
    413, 
    414, 
    415, 
    416, 
    417, 
    418, 
    419, 
    420, 
    421, 
    422, 
    423, 
    424, 
    425, 
    426, 
    427, 
    428, 
    429, 
    430, 
    431, 
    432, 
    433, 
    434, 
    435, 
    436, 
    437, 
    438, 
    439, 
    440, 
    441, 
    442, 
    443, 
    444, 
    445, 
    446, 
    447, 
    448, 
    449, 
    450, 
    451, 
    452, 
    453, 
    454, 
    455, 
    456, 
    457, 
    458, 
    459, 
    460, 
    461, 
    462, 
    463, 
    464, 
    465, 
    466, 
    467, 
    468, 
    469, 
    470, 
    471, 
    472, 
    473, 
    474, 
    475, 
    476, 
    477, 
    478, 
    479, 
    480, 
    481, 
    482, 
    483, 
    484, 
    485, 
    486, 
    487, 
    488, 
    489, 
    490, 
    491, 
    492, 
    493, 
    494, 
    495, 
    496, 
    497, 
    498, 
    499, 
    500, 
    501, 
    502, 
    503, 
    504, 
    505, 
    506, 
    507, 
    508, 
    509, 
    510, 
    511, 
    512, 
    513, 
    514, 
    515, 
    516, 
    517, 
    518, 
    519, 
    520, 
    521, 
    522, 
    523, 
    524, 
    525, 
    526, 
    527, 
    528, 
    529, 
    530, 
    531, 
    532, 
    533, 
    534, 
    535, 
    536, 
    537, 
    538, 
    539, 
    540, 
    541, 
    542, 
    543, 
    544, 
    545, 
    546, 
    547, 
    548, 
    549, 
    550, 
    551, 
    552, 
    553, 
    554, 
    555, 
    556, 
    557, 
    558, 
    559, 
    560, 
    561, 
    562, 
    563, 
    564, 
    565, 
    566, 
    567, 
    568, 
    569, 
    570, 
    571, 
    572, 
    573, 
    574, 
    575, 
    576, 
    577, 
    578, 
    579, 
    580, 
    581, 
    582, 
    583, 
    584, 
    585, 
    586, 
    587, 
    588, 
    589, 
    590, 
    591, 
    592, 
    593, 
    594, 
    595, 
    596, 
    597, 
    598, 
    599, 
    600, 
    601, 
    602, 
    603, 
    604, 
    605, 
    606, 
    607, 
    608, 
    609, 
    610, 
    611, 
    612, 
    613, 
    614, 
    615, 
    616, 
    617, 
    618, 
    619, 
    620, 
    621, 
    622, 
    623, 
    624, 
    625, 
    626, 
    627, 
    628, 
    629, 
    630, 
    631, 
    632, 
    633, 
    634, 
    635, 
    636, 
    637, 
    638, 
    639, 
    640, 
    641, 
    642, 
    643, 
    644, 
    645, 
    646, 
    647, 
    648, 
    649, 
    650, 
    651, 
    652, 
    653, 
    654, 
    655, 
    656, 
    657, 
    658, 
    659, 
    660, 
    661, 
    662, 
    663, 
    664, 
    665, 
    666, 
    667, 
    668, 
    669, 
    670, 
    671, 
    672, 
    673, 
    674, 
    675, 
    676, 
    677, 
    678, 
    679, 
    680, 
    681, 
    682, 
    683, 
    684, 
    685, 
    686, 
    687, 
    688, 
    689, 
    690, 
    691, 
    692, 
    693, 
    694, 
    695, 
    696, 
    697, 
    698, 
    699, 
    700, 
    701, 
    702, 
    703, 
    704, 
    705, 
    706, 
    707, 
    708, 
    709, 
    710, 
    711, 
    712, 
    713, 
    714, 
    715, 
    716, 
    717, 
    718, 
    719, 
    720, 
    721, 
    722, 
    723, 
    724, 
    725, 
    726, 
    727, 
    728, 
    729, 
    730, 
    731, 
    732, 
    733, 
    734, 
    735, 
    736, 
    737, 
    738, 
    739, 
    740, 
    741, 
    742, 
    743, 
    744, 
    745, 
    746, 
    747, 
    748, 
    749, 
    750, 
    751, 
    752, 
    753, 
    754, 
    755, 
    756, 
    757, 
    758, 
    759, 
    760, 
    761, 
    762, 
    763, 
    764, 
    765, 
    766, 
    767, 
    768, 
    769, 
    770, 
    771, 
    772, 
    773, 
    774, 
    775, 
    776, 
    777, 
    778, 
    779, 
    780, 
    781, 
    782, 
    783, 
    784, 
    785, 
    786, 
    787, 
    788, 
    789, 
    790, 
    791, 
    792, 
    793, 
    794, 
    795, 
    796, 
    797, 
    798, 
    799, 
    800, 
    801, 
    802, 
    803, 
    804, 
    805, 
    806, 
    807, 
    808, 
    809, 
    810, 
    811, 
    812, 
    813, 
    814, 
    815, 
    816, 
    817, 
    818, 
    819, 
    820, 
    821, 
    822, 
    823, 
    824, 
    825, 
    826, 
    827, 
    828, 
    829, 
    830, 
    831, 
    832, 
    833, 
    834, 
    835, 
    836, 
    837, 
    838, 
    839, 
    840, 
    841, 
    842, 
    843, 
    844, 
    845, 
    846, 
    847, 
    848, 
    849, 
    850, 
    851, 
    852, 
    853, 
    854, 
    855, 
    856, 
    857, 
    858, 
    859, 
    860, 
    861, 
    862, 
    863, 
    864, 
    865, 
    866, 
    867, 
    868, 
    869, 
    870, 
    871, 
    872, 
    873, 
    874, 
    875, 
    876, 
    877, 
    878, 
    879, 
    880, 
    881, 
    882, 
    883, 
    884, 
    885, 
    886, 
    887, 
    888, 
    889, 
    890, 
    891, 
    892, 
    893, 
    894, 
    895, 
    896, 
    897, 
    898, 
    899, 
    900, 
    901, 
    902, 
    903, 
    904, 
    905, 
    906, 
    907, 
    908, 
    909, 
    910, 
    911, 
    912, 
    913, 
    914, 
    915, 
    916, 
    917, 
    918, 
    919, 
    920, 
    921, 
    922, 
    923, 
    924, 
    925, 
    926, 
    927, 
    928, 
    929, 
    930, 
    931, 
    932, 
    933, 
    934, 
    935, 
    936, 
    937, 
    938, 
    939, 
    940, 
    941, 
    942, 
    943, 
    944, 
    945, 
    946, 
    947, 
    948, 
    949, 
    950, 
    951, 
    952, 
    953, 
    954, 
    955, 
    956, 
    957, 
    958, 
    959, 
    960, 
    961, 
    962, 
    963, 
    964, 
    965, 
    966, 
    967, 
    968, 
    969, 
    970, 
    971, 
    972, 
    973, 
    974, 
    975, 
    976, 
    977, 
    978, 
    979, 
    980, 
    981, 
    982, 
    983, 
    984, 
    985, 
    986, 
    987, 
    988, 
    989, 
    990, 
    991, 
    992, 
    993, 
    994, 
    995, 
    996, 
    997, 
    998, 
    999, 
    1000, 
    1001, 
    1002, 
    1003, 
    1004, 
    1005, 
    1006, 
    1007, 
    1008, 
    1009, 
    1010, 
    1011, 
    1012, 
    1013, 
    1014, 
    1015, 
    1016, 
    1017, 
    1018, 
    1019, 
    1020, 
    1021, 
    1022, 
    1023, 
    1024, 
    1025, 
    1026, 
    1027, 
    1028, 
    1029, 
    1030, 
    1031, 
    1032, 
    1033, 
    1034, 
    1035, 
    1036, 
    1037, 
    1038, 
    1039, 
    1040, 
    1041, 
    1042, 
    1043, 
    1044, 
    1045, 
    1046, 
    1047, 
    1048, 
    1049, 
    1050, 
    1051, 
    1052, 
    1053, 
    1054, 
    1055, 
    1056, 
    1057, 
    1058, 
    1059, 
    1060, 
    1061, 
    1062, 
    1063, 
    1064, 
    1065, 
    1066, 
    1067, 
    1068, 
    1069, 
    1070, 
    1071, 
    1072, 
    1073, 
    1074, 
    1075, 
    1076, 
    1077, 
    1078, 
    1079, 
    1080, 
    1081, 
    1082, 
    1083, 
    1084, 
    1085, 
    1086, 
    1087, 
    1088, 
    1089, 
    1090, 
    1091, 
    1092, 
    1093, 
    1094, 
    1095, 
    1096, 
    1097, 
    1098, 
    1099, 
    1100, 
    1101, 
    1102, 
    1103, 
    1104, 
    1105, 
    1106, 
    1107, 
    1108, 
    1109, 
    1110, 
    1111, 
    1112, 
    1113, 
    1114, 
    1115, 
    1116, 
    1117, 
    1118, 
    1119, 
    1120, 
    1121, 
    1122, 
    1123, 
    1124, 
    1125, 
    1126, 
    1127, 
    1128, 
    1129, 
    1130, 
    1131, 
    1132, 
    1133, 
    1134, 
    1135, 
    1136, 
    1137, 
    1138, 
    1139, 
    1140, 
    1141, 
    1142, 
    1143, 
    1144, 
    1145, 
    1146, 
    1147, 
    1148, 
    1149, 
    1150, 
    1151, 
    1152, 
    1153, 
    1154, 
    1155, 
    1156, 
    1157, 
    1158, 
    1159, 
    1160, 
    1161, 
    1162, 
    1163, 
    1164, 
    1165, 
    1166, 
    1167, 
    1168, 
    1169, 
    1170, 
    1171, 
    1172, 
    1173, 
    1174, 
    1175, 
    1176, 
    1177, 
    1178, 
    1179, 
    1180, 
    1181, 
    1182, 
    1183, 
    1184, 
    1185, 
    1186, 
    1187, 
    1188, 
    1189, 
    1190, 
    1191, 
    1192, 
    1193, 
    1194, 
    1195, 
    1196, 
    1197, 
    1198, 
    1199, 
    1200, 
    1201, 
    1202, 
    1203, 
    1204, 
    1205, 
    1206, 
    1207, 
    1208, 
    1209, 
    1210, 
    1211, 
    1212, 
    1213, 
    1214, 
    1215, 
    1216, 
    1217, 
    1218, 
    1219, 
    1220, 
    1221, 
    1222, 
    1223, 
    1224, 
    1225, 
    1226, 
    1227, 
    1228, 
    1229, 
    1230, 
    1231, 
    1232, 
    1233, 
    1234, 
    1235, 
    1236, 
    1237, 
    1238, 
    1239, 
    1240, 
    1241, 
    1242, 
    1243, 
    1244, 
    1245, 
    1246, 
    1247, 
    1248, 
    1249, 
    1250, 
    1251, 
    1252, 
    1253, 
    1254, 
    1255, 
    1256, 
    1257, 
    1258, 
    1259, 
    1260, 
    1261, 
    1262, 
    1263, 
    1264, 
    1265, 
    1266, 
    1267, 
    1268, 
    1269, 
    1270, 
    1271, 
    1272, 
    1273, 
    1274, 
    1275, 
    1276, 
    1277, 
    1278, 
    1279, 
    1280, 
    1281, 
    1282, 
    1283, 
    1284, 
    1285, 
    1286, 
    1287, 
    1288, 
    1289, 
    1290, 
    1291, 
    1292, 
    1293, 
    1294, 
    1295, 
    1296, 
    1297, 
    1298, 
    1299, 
    1300, 
    1301, 
    1302, 
    1303, 
    1304, 
    1305, 
    1306, 
    1307, 
    1308, 
    1309, 
    1310, 
    1311, 
    1312, 
    1313, 
    1314, 
    1315, 
    1316, 
    1317, 
    1318, 
    1319, 
    1320, 
    1321, 
    1322, 
    1323, 
    1324, 
    1325, 
    1326, 
    1327, 
    1328, 
    1329, 
    1330, 
    1331, 
    1332, 
    1333, 
    1334, 
    1335, 
    1336, 
    1337, 
    1338, 
    1339, 
    1340, 
    1341, 
    1342, 
    1343, 
    1344, 
    1345, 
    1346, 
    1347, 
    1348, 
    1349, 
    1350, 
    1351, 
    1352, 
    1353, 
    1354, 
    1355, 
    1356, 
    1357, 
    1358, 
    1359, 
    1360, 
    1361, 
    1362, 
    1363, 
    1364, 
    1365, 
    1366, 
    1367, 
    1368, 
    1369, 
    1370, 
    1371, 
    1372, 
    1373, 
    1374, 
    1375, 
    1376, 
    1377, 
    1378, 
    1379, 
    1380, 
    1381, 
    1382, 
    1383, 
    1384, 
    1385, 
    1386, 
    1387, 
    1388, 
    1389, 
    1390, 
    1391, 
    1392, 
    1393, 
    1394, 
    1395, 
    1396, 
    1397, 
    1398, 
    1399, 
    1400, 
    1401, 
    1402, 
    1403, 
    1404, 
    1405, 
    1406, 
    1407, 
    1408, 
    1409, 
    1410, 
    1411, 
    1412, 
    1413, 
    1414, 
    1415, 
    1416, 
    1417, 
    1418, 
    1419, 
    1420, 
    1421, 
    1422, 
    1423, 
    1424, 
    1425, 
    1426, 
    1427, 
    1428, 
    1429, 
    1430, 
    1431, 
    1432, 
    1433, 
    1434, 
    1435, 
    1436, 
    1437, 
    1438, 
    1439, 
    1440, 
    1441, 
    1442, 
    1443, 
    1444, 
    1445, 
    1446, 
    1447, 
    1448, 
    1449, 
    1450, 
    1451, 
    1452, 
    1453, 
    1454, 
    1455, 
    1456, 
    1457, 
    1458, 
    1459, 
    1460, 
    1461, 
    1462, 
    1463, 
    1464, 
    1465, 
    1466, 
    1467, 
    1468, 
    1469, 
    1470, 
    1471, 
    1472, 
    1473, 
    1474, 
    1475, 
    1476, 
    1477, 
    1478, 
    1479, 
    1480, 
    1481, 
    1482, 
    1483, 
    1484, 
    1485, 
    1486, 
    1487, 
    1488, 
    1489, 
    1490, 
    1491, 
    1492, 
    1493, 
    1494, 
    1495, 
    1496, 
    1497, 
    1498, 
    1499, 
    1500, 
    1501, 
    1502, 
    1503, 
    1504, 
    1505, 
    1506, 
    1507, 
    1508, 
    1509, 
    1510, 
    1511, 
    1512, 
    1513, 
    1514, 
    1515, 
    1516, 
    1517, 
    1518, 
    1519, 
    1520, 
    1521, 
    1522, 
    1523, 
    1524, 
    1525, 
    1526, 
    1527, 
    1528, 
    1529, 
    1530, 
    1531, 
    1532, 
    1533, 
    1534, 
    1535, 
    1536, 
    1537, 
    1538, 
    1539, 
    1540, 
    1541, 
    1542, 
    1543, 
    1544, 
    1545, 
    1546, 
    1547, 
    1548, 
    1549, 
    1550, 
    1551, 
    1552, 
    1553, 
    1554, 
    1555, 
    1556, 
    1557, 
    1558, 
    1559, 
    1560, 
    1561, 
    1562, 
    1563, 
    1564, 
    1565, 
    1566, 
    1567, 
    1568, 
    1569, 
    1570, 
    1571, 
    1572, 
    1573, 
    1574, 
    1575, 
    1576, 
    1577, 
    1578, 
    1579, 
    1580, 
    1581, 
    1582, 
    1583, 
    1584, 
    1585, 
    1586, 
    1587, 
    1588, 
    1589, 
    1590, 
    1591, 
    1592, 
    1593, 
    1594, 
    1595, 
    1596, 
    1597, 
    1598, 
    1599, 
    1600, 
    1601, 
    1602, 
    1603, 
    1604, 
    1605, 
    1606, 
    1607, 
    1608, 
    1609, 
    1610, 
    1611, 
    1612, 
    1613, 
    1614, 
    1615, 
    1616, 
    1617, 
    1618, 
    1619, 
    1620, 
    1621, 
    1622, 
    1623, 
    1624, 
    1625, 
    1626, 
    1627, 
    1628, 
    1629, 
    1630, 
    1631, 
    1632, 
    1633, 
    1634, 
    1635, 
    1636, 
    1637, 
    1638, 
    1639, 
    1640, 
    1641, 
    1642, 
    1643, 
    1644, 
    1645, 
    1646, 
    1647, 
    1648, 
    1649, 
    1650, 
    1651, 
    1652, 
    1653, 
    1654, 
    1655, 
    1656, 
    1657, 
    1658, 
    1659, 
    1660, 
    1661, 
    1662, 
    1663, 
    1664, 
    1665, 
    1666, 
    1667, 
    1668, 
    1669, 
    1670, 
    1671, 
    1672, 
    1673, 
    1674, 
    1675, 
    1676, 
    1677, 
    1678, 
    1679, 
    1680, 
    1681, 
    1682, 
    1683, 
    1684, 
    1685, 
    1686, 
    1687, 
    1688, 
    1689, 
    1690, 
    1691, 
    1692, 
    1693, 
    1694, 
    1695, 
    1696, 
    1697, 
    1698, 
    1699, 
    1700, 
    1701, 
    1702, 
    1703, 
    1704, 
    1705, 
    1706, 
    1707, 
    1708, 
    1709, 
    1710, 
    1711, 
    1712, 
    1713, 
    1714, 
    1715, 
    1716, 
    1717, 
    1718, 
    1719, 
    1720, 
    1721, 
    1722, 
    1723, 
    1724, 
    1725, 
    1726, 
    1727, 
    1728, 
    1729, 
    1730, 
    1731, 
    1732, 
    1733, 
    1734, 
    1735, 
    1736, 
    1737, 
    1738, 
    1739, 
    1740, 
    1741, 
    1742, 
    1743, 
    1744, 
    1745, 
    1746, 
    1747, 
    1748, 
    1749, 
    1750, 
    1751, 
    1752, 
    1753, 
    1754, 
    1755, 
    1756, 
    1757, 
    1758, 
    1759, 
    1760, 
    1761, 
    1762, 
    1763, 
    1764, 
    1765, 
    1766, 
    1767, 
    1768, 
    1769, 
    1770, 
    1771, 
    1772, 
    1773, 
    1774, 
    1775, 
    1776, 
    1777, 
    1778, 
    1779, 
    1780, 
    1781, 
    1782, 
    1783, 
    1784, 
    1785, 
    1786, 
    1787, 
    1788, 
    1789, 
    1790, 
    1791, 
    1792, 
    1793, 
    1794, 
    1795, 
    1796, 
    1797, 
    1798, 
    1799, 
    1800, 
    1801, 
    1802, 
    1803, 
    1804, 
    1805, 
    1806, 
    1807, 
    1808, 
    1809, 
    1810, 
    1811, 
    1812, 
    1813, 
    1814, 
    1815, 
    1816, 
    1817, 
    1818, 
    1819, 
    1820, 
    1821, 
    1822, 
    1823, 
    1824, 
    1825, 
    1826, 
    1827, 
    1828, 
    1829, 
    1830, 
    1831, 
    1832, 
    1833, 
    1834, 
    1835, 
    1836, 
    1837, 
    1838, 
    1839, 
    1840, 
    1841, 
    1842, 
    1843, 
    1844, 
    1845, 
    1846, 
    1847, 
    1848, 
    1849, 
    1850, 
    1851, 
    1852, 
    1853, 
    1854, 
    1855, 
    1856, 
    1857, 
    1858, 
    1859, 
    1860, 
    1861, 
    1862, 
    1863, 
    1864, 
    1865, 
    1866, 
    1867, 
    1868, 
    1869, 
    1870, 
    1871, 
    1872, 
    1873, 
    1874, 
    1875, 
    1876, 
    1877, 
    1878, 
    1879, 
    1880, 
    1881, 
    1882, 
    1883, 
    1884, 
    1885, 
    1886, 
    1887, 
    1888, 
    1889, 
    1890, 
    1891, 
    1892, 
    1893, 
    1894, 
    1895, 
    1896, 
    1897, 
    1898, 
    1899, 
    1900, 
    1901, 
    1902, 
    1903, 
    1904, 
    1905, 
    1906, 
    1907, 
    1908, 
    1909, 
    1910, 
    1911, 
    1912, 
    1913, 
    1914, 
    1915, 
    1916, 
    1917, 
    1918, 
    1919, 
    1920, 
    1921, 
    1922, 
    1923, 
    1924, 
    1925, 
    1926, 
    1927, 
    1928, 
    1929, 
    1930, 
    1931, 
    1932, 
    1933, 
    1934, 
    1935, 
    1936, 
    1937, 
    1938, 
    1939, 
    1940, 
    1941, 
    1942, 
    1943, 
    1944, 
    1945, 
    1946, 
    1947, 
    1948, 
    1949, 
    1950, 
    1951, 
    1952, 
    1953, 
    1954, 
    1955, 
    1956, 
    1957, 
    1958, 
    1959, 
    1960, 
    1961, 
    1962, 
    1963, 
    1964, 
    1965, 
    1966, 
    1967, 
    1968, 
    1969, 
    1970, 
    1971, 
    1972, 
    1973, 
    1974, 
    1975, 
    1976, 
    1977, 
    1978, 
    1979, 
    1980, 
    1981, 
    1982, 
    1983, 
    1984, 
    1985, 
    1986, 
    1987, 
    1988, 
    1989, 
    1990, 
    1991, 
    1992, 
    1993, 
    1994, 
    1995, 
    1996, 
    1997, 
    1998, 
    1999, 
    2000, 
    2001, 
    2002, 
    2003, 
    2004, 
    2005, 
    2006, 
    2007, 
    2008, 
    2009, 
    2010, 
    2011, 
    2012, 
    2013, 
    2014, 
    2015, 
    2016, 
    2017, 
    2018, 
    2019, 
    2020, 
    2021, 
    2022, 
    2023, 
    2024, 
    2025, 
    2026, 
    2027, 
    2028, 
    2029, 
    2030, 
    2031, 
    2032, 
    2033, 
    2034, 
    2035, 
    2036, 
    2037, 
    2038, 
    2039, 
    2040, 
    2041, 
    2042, 
    2043, 
    2044, 
    2045, 
    2046, 
    2047, 
    2048, 
    2049, 
    2050, 
    2051, 
    2052, 
    2053, 
    2054, 
    2055, 
    2056, 
    2057, 
    2058, 
    2059, 
    2060, 
    2061, 
    2062, 
    2063, 
    2064, 
    2065, 
    2066, 
    2067, 
    2068, 
    2069, 
    2070, 
    2071, 
    2072, 
    2073, 
    2074, 
    2075, 
    2076, 
    2077, 
    2078, 
    2079, 
    2080, 
    2081, 
    2082, 
    2083, 
    2084, 
    2085, 
    2086, 
    2087, 
    2088, 
    2089, 
    2090, 
    2091, 
    2092, 
    2093, 
    2094, 
    2095, 
    2096, 
    2097, 
    2098, 
    2099, 
    2100, 
    2101, 
    2102, 
    2103, 
    2104, 
    2105, 
    2106, 
    2107, 
    2108, 
    2109, 
    2110, 
    2111, 
    2112, 
    2113, 
    2114, 
    2115, 
    2116, 
    2117, 
    2118, 
    2119, 
    2120, 
    2121, 
    2122, 
    2123, 
    2124, 
    2125, 
    2126, 
    2127, 
    2128, 
    2129, 
    2130, 
    2131, 
    2132, 
    2133, 
    2134, 
    2135, 
    2136, 
    2137, 
    2138, 
    2139, 
    2140, 
    2141, 
    2142, 
    2143, 
    2144, 
    2145, 
    2146, 
    2147, 
    2148, 
    2149, 
    2150, 
    2151, 
    2152, 
    2153, 
    2154, 
    2155, 
    2156, 
    2157, 
    2158, 
    2159, 
    2160, 
    2161, 
    2162, 
    2163, 
    2164, 
    2165, 
    2166, 
    2167, 
    2168, 
    2169, 
    2170, 
    2171, 
    2172, 
    2173, 
    2174, 
    2175, 
    2176, 
    2177, 
    2178, 
    2179, 
    2180, 
    2181, 
    2182, 
    2183, 
    2184, 
    2185, 
    2186, 
    2187, 
    2188, 
    2189, 
    2190, 
    2191, 
    2192, 
    2193, 
    2194, 
    2195, 
    2196, 
    2197, 
    2198, 
    2199, 
    2200, 
    2201, 
    2202, 
    2203, 
    2204, 
    2205, 
    2206, 
    2207, 
    2208, 
    2209, 
    2210, 
    2211, 
    2212, 
    2213, 
    2214, 
    2215, 
    2216, 
    2217, 
    2218, 
    2219, 
    2220, 
    2221, 
    2222, 
    2223, 
    2224, 
    2225, 
    2226, 
    2227, 
    2228, 
    2229, 
    2230, 
    2231, 
    2232, 
    2233, 
    2234, 
    2235, 
    2236, 
    2237, 
    2238, 
    2239, 
    2240, 
    2241, 
    2242, 
    2243, 
    2244, 
    2245, 
    2246, 
    2247, 
    2248, 
    2249, 
    2250, 
    2251, 
    2252, 
    2253, 
    2254, 
    2255, 
    2256, 
    2257, 
    2258, 
    2259, 
    2260, 
    2261, 
    2262, 
    2263, 
    2264, 
    2265, 
    2266, 
    2267, 
    2268, 
    2269, 
    2270, 
    2271, 
    2272, 
    2273, 
    2274, 
    2275, 
    2276, 
    2277, 
    2278, 
    2279, 
    2280, 
    2281, 
    2282, 
    2283, 
    2284, 
    2285, 
    2286, 
    2287, 
    2288, 
    2289, 
    2290, 
    2291, 
    2292, 
    2293, 
    2294, 
    2295, 
    2296, 
    2297, 
    2298, 
    2299, 
    2300, 
    2301, 
    2302, 
    2303, 
    2304, 
    2305, 
    2306, 
    2307, 
    2308, 
    2309, 
    2310, 
    2311, 
    2312, 
    2313, 
    2314, 
    2315, 
    2316, 
    2317, 
    2318, 
    2319, 
    2320, 
    2321, 
    2322, 
    2323, 
    2324, 
    2325, 
    2326, 
    2327, 
    2328, 
    2329, 
    2330, 
    2331, 
    2332, 
    2333, 
    2334, 
    2335, 
    2336, 
    2337, 
    2338, 
    2339, 
    2340, 
    2341, 
    2342, 
    2343, 
    2344, 
    2345, 
    2346, 
    2347, 
    2348, 
    2349, 
    2350, 
    2351, 
    2352, 
    2353, 
    2354, 
    2355, 
    2356, 
    2357, 
    2358, 
    2359, 
    2360, 
    2361, 
    2362, 
    2363, 
    2364, 
    2365, 
    2366, 
    2367, 
    2368, 
    2369, 
    2370, 
    2371, 
    2372, 
    2373, 
    2374, 
    2375, 
    2376, 
    2377, 
    2378, 
    2379, 
    2380, 
    2381, 
    2382, 
    2383, 
    2384, 
    2385, 
    2386, 
    2387, 
    2388, 
    2389, 
    2390, 
    2391, 
    2392, 
    2393, 
    2394, 
    2395, 
    2396, 
    2397, 
    2398, 
    2399, 
    2400, 
    2401, 
    2402, 
    2403, 
    2404, 
    2405, 
    2406, 
    2407, 
    2408, 
    2409, 
    2410, 
    2411, 
    2412, 
    2413, 
    2414, 
    2415, 
    2416, 
    2417, 
    2418, 
    2419, 
    2420, 
    2421, 
    2422, 
    2423, 
    2424, 
    2425, 
    2426, 
    2427, 
    2428, 
    2429, 
    2430, 
    2431, 
    2432, 
    2433, 
    2434, 
    2435, 
    2436, 
    2437, 
    2438, 
    2439, 
    2440, 
    2441, 
    2442, 
    2443, 
    2444, 
    2445, 
    2446, 
    2447, 
    2448, 
    2449, 
    2450, 
    2451, 
    2452, 
    2453, 
    2454, 
    2455, 
    2456, 
    2457, 
    2458, 
    2459, 
    2460, 
    2461, 
    2462, 
    2463, 
    2464, 
    2465, 
    2466, 
    2467, 
    2468, 
    2469, 
    2470, 
    2471, 
    2472, 
    2473, 
    2474, 
    2475, 
    2476, 
    2477, 
    2478, 
    2479, 
    2480, 
    2481, 
    2482, 
    2483, 
    2484, 
    2485, 
    2486, 
    2487, 
    2488, 
    2489, 
    2490, 
    2491, 
    2492, 
    2493, 
    2494, 
    2495, 
    2496, 
    2497, 
    2498, 
    2499, 
    2500, 
    2501, 
    2502, 
    2503, 
    2504, 
    2505, 
    2506, 
    2507, 
    2508, 
    2509, 
    2510, 
    2511, 
    2512, 
    2513, 
    2514, 
    2515, 
    2516, 
    2517, 
    2518, 
    2519, 
    2520, 
    2521, 
    2522, 
    2523, 
    2524, 
    2525, 
    2526, 
    2527, 
    2528, 
    2529, 
    2530, 
    2531, 
    2532, 
    2533, 
    2534, 
    2535, 
    2536, 
    2537, 
    2538, 
    2539, 
    2540, 
    2541, 
    2542, 
    2543, 
    2544, 
    2545, 
    2546, 
    2547, 
    2548, 
    2549, 
    2550, 
    2551, 
    2552, 
    2553, 
    2554, 
    2555, 
    2556, 
    2557, 
    2558, 
    2559, 
    2560, 
    2561, 
    2562, 
    2563, 
    2564, 
    2565, 
    2566, 
    2567, 
    2568, 
    2569, 
    2570, 
    2571, 
    2572, 
    2573, 
    2574, 
    2575, 
    2576, 
    2577, 
    2578, 
    2579, 
    2580, 
    2581, 
    2582, 
    2583, 
    2584, 
    2585, 
    2586, 
    2587, 
    2588, 
    2589, 
    2590, 
    2591, 
    2592, 
    2593, 
    2594, 
    2595, 
    2596, 
    2597, 
    2598, 
    2599, 
    2600, 
    2601, 
    2602, 
    2603, 
    2604, 
    2605, 
    2606, 
    2607, 
    2608, 
    2609, 
    2610, 
    2611, 
    2612, 
    2613, 
    2614, 
    2615, 
    2616, 
    2617, 
    2618, 
    2619, 
    2620, 
    2621, 
    2622, 
    2623, 
    2624, 
    2625, 
    2626, 
    2627, 
    2628, 
    2629, 
    2630, 
    2631, 
    2632, 
    2633, 
    2634, 
    2635, 
    2636, 
    2637, 
    2638, 
    2639, 
    2640, 
    2641, 
    2642, 
    2643, 
    2644, 
    2645, 
    2646, 
    2647, 
    2648, 
    2649, 
    2650, 
    2651, 
    2652, 
    2653, 
    2654, 
    2655, 
    2656, 
    2657, 
    2658, 
    2659, 
    2660, 
    2661, 
    2662, 
    2663, 
    2664, 
    2665, 
    2666, 
    2667, 
    2668, 
    2669, 
    2670, 
    2671, 
    2672, 
    2673, 
    2674, 
    2675, 
    2676, 
    2677, 
    2678, 
    2679, 
    2680, 
    2681, 
    2682, 
    2683, 
    2684, 
    2685, 
    2686, 
    2687, 
    2688, 
    2689, 
    2690, 
    2691, 
    2692, 
    2693, 
    2694, 
    2695, 
    2696, 
    2697, 
    2698, 
    2699, 
    2700, 
    2701, 
    2702, 
    2703, 
    2704, 
    2705, 
    2706, 
    2707, 
    2708, 
    2709, 
    2710, 
    2711, 
    2712, 
    2713, 
    2714, 
    2715, 
    2716, 
    2717, 
    2718, 
    2719, 
    2720, 
    2721, 
    2722, 
    2723, 
    2724, 
    2725, 
    2726, 
    2727, 
    2728, 
    2729, 
    2730, 
    2731, 
    2732, 
    2733, 
    2734, 
    2735, 
    2736, 
    2737, 
    2738, 
    2739, 
    2740, 
    2741, 
    2742, 
    2743, 
    2744, 
    2745, 
    2746, 
    2747, 
    2748, 
    2749, 
    2750, 
    2751, 
    2752, 
    2753, 
    2754, 
    2755, 
    2756, 
    2757, 
    2758, 
    2759, 
    2760, 
    2761, 
    2762, 
    2763, 
    2764, 
    2765, 
    2766, 
    2767, 
    2768, 
    2769, 
    2770, 
    2771, 
    2772, 
    2773, 
    2774, 
    2775, 
    2776, 
    2777, 
    2778, 
    2779, 
    2780, 
    2781, 
    2782, 
    2783, 
    2784, 
    2785, 
    2786, 
    2787, 
    2788, 
    2789, 
    2790, 
    2791, 
    2792, 
    2793, 
    2794, 
    2795, 
    2796, 
    2797, 
    2798, 
    2799, 
    2800, 
    2801, 
    2802, 
    2803, 
    2804, 
    2805, 
    2806, 
    2807, 
    2808, 
    2809, 
    2810, 
    2811, 
    2812, 
    2813, 
    2814, 
    2815, 
    2816, 
    2817, 
    2818, 
    2819, 
    2820, 
    2821, 
    2822, 
    2823, 
    2824, 
    2825, 
    2826, 
    2827, 
    2828, 
    2829, 
    2830, 
    2831, 
    2832, 
    2833, 
    2834, 
    2835, 
    2836, 
    2837, 
    2838, 
    2839, 
    2840, 
    2841, 
    2842, 
    2843, 
    2844, 
    2845, 
    2846, 
    2847, 
    2848, 
    2849, 
    2850, 
    2851, 
    2852, 
    2853, 
    2854, 
    2855, 
    2856, 
    2857, 
    2858, 
    2859, 
    2860, 
    2861, 
    2862, 
    2863, 
    2864, 
    2865, 
    2866, 
    2867, 
    2868, 
    2869, 
    2870, 
    2871, 
    2872, 
    2873, 
    2874, 
    2875, 
    2876, 
    2877, 
    2878, 
    2879, 
    2880, 
    2881, 
    2882, 
    2883, 
    2884, 
    2885, 
    2886, 
    2887, 
    2888, 
    2889, 
    2890, 
    2891, 
    2892, 
    2893, 
    2894, 
    2895, 
    2896, 
    2897, 
    2898, 
    2899, 
    2900, 
    2901, 
    2902, 
    2903, 
    2904, 
    2905, 
    2906, 
    2907, 
    2908, 
    2909, 
    2910, 
    2911, 
    2912, 
    2913, 
    2914, 
    2915, 
    2916, 
    2917, 
    2918, 
    2919, 
    2920, 
    2921, 
    2922, 
    2923, 
    2924, 
    2925, 
    2926, 
    2927, 
    2928, 
    2929, 
    2930, 
    2931, 
    2932, 
    2933, 
    2934, 
    2935, 
    2936, 
    2937, 
    2938, 
    2939, 
    2940, 
    2941, 
    2942, 
    2943, 
    2944, 
    2945, 
    2946, 
    2947, 
    2948, 
    2949, 
    2950, 
    2951, 
    2952, 
    2953, 
    2954, 
    2955, 
    2956, 
    2957, 
    2958, 
    2959, 
    2960, 
    2961, 
    2962, 
    2963, 
    2964, 
    2965, 
    2966, 
    2967, 
    2968, 
    2969, 
    2970, 
    2971, 
    2972, 
    2973, 
    2974, 
    2975, 
    2976, 
    2977, 
    2978, 
    2979, 
    2980, 
    2981, 
    2982, 
    2983, 
    2984, 
    2985, 
    2986, 
    2987, 
    2988, 
    2989, 
    2990, 
    2991, 
    2992, 
    2993, 
    2994, 
    2995, 
    2996, 
    2997, 
    2998, 
    2999, 
    3000, 
    3001, 
    3002, 
    3003, 
    3004, 
    3005, 
    3006, 
    3007, 
    3008, 
    3009, 
    3010, 
    3011, 
    3012, 
    3013, 
    3014, 
    3015, 
    3016, 
    3017, 
    3018, 
    3019, 
    3020, 
    3021, 
    3022, 
    3023, 
    3024, 
    3025, 
    3026, 
    3027, 
    3028, 
    3029, 
    3030, 
    3031, 
    3032, 
    3033, 
    3034, 
    3035, 
    3036, 
    3037, 
    3038, 
    3039, 
    3040, 
    3041, 
    3042, 
    3043, 
    3044, 
    3045, 
    3046, 
    3047, 
    3048, 
    3049, 
    3050, 
    3051, 
    3052, 
    3053, 
    3054, 
    3055, 
    3056, 
    3057, 
    3058, 
    3059, 
    3060, 
    3061, 
    3062, 
    3063, 
    3064, 
    3065, 
    3066, 
    3067, 
    3068, 
    3069, 
    3070, 
    3071, 
    3072, 
    3073, 
    3074, 
    3075, 
    3076, 
    3077, 
    3078, 
    3079, 
    3080, 
    3081, 
    3082, 
    3083, 
    3084, 
    3085, 
    3086, 
    3087, 
    3088, 
    3089, 
    3090, 
    3091, 
    3092, 
    3093, 
    3094, 
    3095, 
    3096, 
    3097, 
    3098, 
    3099, 
    3100, 
    3101, 
    3102, 
    3103, 
    3104, 
    3105, 
    3106, 
    3107, 
    3108, 
    3109, 
    3110, 
    3111, 
    3112, 
    3113, 
    3114, 
    3115, 
    3116, 
    3117, 
    3118, 
    3119, 
    3120, 
    3121, 
    3122, 
    3123, 
    3124, 
    3125, 
    3126, 
    3127, 
    3128, 
    3129, 
    3130, 
    3131, 
    3132, 
    3133, 
    3134, 
    3135, 
    3136, 
    3137, 
    3138, 
    3139, 
    3140, 
    3141, 
    3142, 
    3143, 
    3144, 
    3145, 
    3146, 
    3147, 
    3148, 
    3149, 
    3150, 
    3151, 
    3152, 
    3153, 
    3154, 
    3155, 
    3156, 
    3157, 
    3158, 
    3159, 
    3160, 
    3161, 
    3162, 
    3163, 
    3164, 
    3165, 
    3166, 
    3167, 
    3168, 
    3169, 
    3170, 
    3171, 
    3172, 
    3173, 
    3174, 
    3175, 
    3176, 
    3177, 
    3178, 
    3179, 
    3180, 
    3181, 
    3182, 
    3183, 
    3184, 
    3185, 
    3186, 
    3187, 
    3188, 
    3189, 
    3190, 
    3191, 
    3192, 
    3193, 
    3194, 
    3195, 
    3196, 
    3197, 
    3198, 
    3199, 
    3200, 
    3201, 
    3202, 
    3203, 
    3204, 
    3205, 
    3206, 
    3207, 
    3208, 
    3209, 
    3210, 
    3211, 
    3212, 
    3213, 
    3214, 
    3215, 
    3216, 
    3217, 
    3218, 
    3219, 
    3220, 
    3221, 
    3222, 
    3223, 
    3224, 
    3225, 
    3226, 
    3227, 
    3228, 
    3229, 
    3230, 
    3231, 
    3232, 
    3233, 
    3234, 
    3235, 
    3236, 
    3237, 
    3238, 
    3239, 
    3240, 
    3241, 
    3242, 
    3243, 
    3244, 
    3245, 
    3246, 
    3247, 
    3248, 
    3249, 
    3250, 
    3251, 
    3252, 
    3253, 
    3254, 
    3255, 
    3256, 
    3257, 
    3258, 
    3259, 
    3260, 
    3261, 
    3262, 
    3263, 
    3264, 
    3265, 
    3266, 
    3267, 
    3268, 
    3269, 
    3270, 
    3271, 
    3272, 
    3273, 
    3274, 
    3275, 
    3276, 
    3277, 
    3278, 
    3279, 
    3280, 
    3281, 
    3282, 
    3283, 
    3284, 
    3285, 
    3286, 
    3287, 
    3288, 
    3289, 
    3290, 
    3291, 
    3292, 
    3293, 
    3294, 
    3295, 
    3296, 
    3297, 
    3298, 
    3299, 
    3300, 
    3301, 
    3302, 
    3303, 
    3304, 
    3305, 
    3306, 
    3307, 
    3308, 
    3309, 
    3310, 
    3311, 
    3312, 
    3313, 
    3314, 
    3315, 
    3316, 
    3317, 
    3318, 
    3319, 
    3320, 
    3321, 
    3322, 
    3323, 
    3324, 
    3325, 
    3326, 
    3327, 
    3328, 
    3329, 
    3330, 
    3331, 
    3332, 
    3333, 
    3334, 
    3335, 
    3336, 
    3337, 
    3338, 
    3339, 
    3340, 
    3341, 
    3342, 
    3343, 
    3344, 
    3345, 
    3346, 
    3347, 
    3348, 
    3349, 
    3350, 
    3351, 
    3352, 
    3353, 
    3354, 
    3355, 
    3356, 
    3357, 
    3358, 
    3359, 
    3360, 
    3361, 
    3362, 
    3363, 
    3364, 
    3365, 
    3366, 
    3367, 
    3368, 
    3369, 
    3370, 
    3371, 
    3372, 
    3373, 
    3374, 
    3375, 
    3376, 
    3377, 
    3378, 
    3379, 
    3380, 
    3381, 
    3382, 
    3383, 
    3384, 
    3385, 
    3386, 
    3387, 
    3388, 
    3389, 
    3390, 
    3391, 
    3392, 
    3393, 
    3394, 
    3395, 
    3396, 
    3397, 
    3398, 
    3399, 
    3400, 
    3401, 
    3402, 
    3403, 
    3404, 
    3405, 
    3406, 
    3407, 
    3408, 
    3409, 
    3410, 
    3411, 
    3412, 
    3413, 
    3414, 
    3415, 
    3416, 
    3417, 
    3418, 
    3419, 
    3420, 
    3421, 
    3422, 
    3423, 
    3424, 
    3425, 
    3426, 
    3427, 
    3428, 
    3429, 
    3430, 
    3431, 
    3432, 
    3433, 
    3434, 
    3435, 
    3436, 
    3437, 
    3438, 
    3439, 
    3440, 
    3441, 
    3442, 
    3443, 
    3444, 
    3445, 
    3446, 
    3447, 
    3448, 
    3449, 
    3450, 
    3451, 
    3452, 
    3453, 
    3454, 
    3455, 
    3456, 
    3457, 
    3458, 
    3459, 
    3460, 
    3461, 
    3462, 
    3463, 
    3464, 
    3465, 
    3466, 
    3467, 
    3468, 
    3469, 
    3470, 
    3471, 
    3472, 
    3473, 
    3474, 
    3475, 
    3476, 
    3477, 
    3478, 
    3479, 
    3480, 
    3481, 
    3482, 
    3483, 
    3484, 
    3485, 
    3486, 
    3487, 
    3488, 
    3489, 
    3490, 
    3491, 
    3492, 
    3493, 
    3494, 
    3495, 
    3496, 
    3497, 
    3498, 
    3499, 
    3500, 
    3501, 
    3502, 
    3503, 
    3504, 
    3505, 
    3506, 
    3507, 
    3508, 
    3509, 
    3510, 
    3511, 
    3512, 
    3513, 
    3514, 
    3515, 
    3516, 
    3517, 
    3518, 
    3519, 
    3520, 
    3521, 
    3522, 
    3523, 
    3524, 
    3525, 
    3526, 
    3527, 
    3528, 
    3529, 
    3530, 
    3531, 
    3532, 
    3533, 
    3534, 
    3535, 
    3536, 
    3537, 
    3538, 
    3539, 
    3540, 
    3541, 
    3542, 
    3543, 
    3544, 
    3545, 
    3546, 
    3547, 
    3548, 
    3549, 
    3550, 
    3551, 
    3552, 
    3553, 
    3554, 
    3555, 
    3556, 
    3557, 
    3558, 
    3559, 
    3560, 
    3561, 
    3562, 
    3563, 
    3564, 
    3565, 
    3566, 
    3567, 
    3568, 
    3569, 
    3570, 
    3571, 
    3572, 
    3573, 
    3574, 
    3575, 
    3576, 
    3577, 
    3578, 
    3579, 
    3580, 
    3581, 
    3582, 
    3583, 
    3584, 
    3585, 
    3586, 
    3587, 
    3588, 
    3589, 
    3590, 
    3591, 
    3592, 
    3593, 
    3594, 
    3595, 
    3596, 
    3597, 
    3598, 
    3599, 
    3600, 
    3601, 
    3602, 
    3603, 
    3604, 
    3605, 
    3606, 
    3607, 
    3608, 
    3609, 
    3610, 
    3611, 
    3612, 
    3613, 
    3614, 
    3615, 
    3616, 
    3617, 
    3618, 
    3619, 
    3620, 
    3621, 
    3622, 
    3623, 
    3624, 
    3625, 
    3626, 
    3627, 
    3628, 
    3629, 
    3630, 
    3631, 
    3632, 
    3633, 
    3634, 
    3635, 
    3636, 
    3637, 
    3638, 
    3639, 
    3640, 
    3641, 
    3642, 
    3643, 
    3644, 
    3645, 
    3646, 
    3647, 
    3648, 
    3649, 
    3650, 
    3651, 
    3652, 
    3653, 
    3654, 
    3655, 
    3656, 
    3657, 
    3658, 
    3659, 
    3660, 
    3661, 
    3662, 
    3663, 
    3664, 
    3665, 
    3666, 
    3667, 
    3668, 
    3669, 
    3670, 
    3671, 
    3672, 
    3673, 
    3674, 
    3675, 
    3676, 
    3677, 
    3678, 
    3679, 
    3680, 
    3681, 
    3682, 
    3683, 
    3684, 
    3685, 
    3686, 
    3687, 
    3688, 
    3689, 
    3690, 
    3691, 
    3692, 
    3693, 
    3694, 
    3695, 
    3696, 
    3697, 
    3698, 
    3699, 
    3700, 
    3701, 
    3702, 
    3703, 
    3704, 
    3705, 
    3706, 
    3707, 
    3708, 
    3709, 
    3710, 
    3711, 
    3712, 
    3713, 
    3714, 
    3715, 
    3716, 
    3717, 
    3718, 
    3719, 
    3720, 
    3721, 
    3722, 
    3723, 
    3724, 
    3725, 
    3726, 
    3727, 
    3728, 
    3729, 
    3730, 
    3731, 
    3732, 
    3733, 
    3734, 
    3735, 
    3736, 
    3737, 
    3738, 
    3739, 
    3740, 
    3741, 
    3742, 
    3743, 
    3744, 
    3745, 
    3746, 
    3747, 
    3748, 
    3749, 
    3750, 
    3751, 
    3752, 
    3753, 
    3754, 
    3755, 
    3756, 
    3757, 
    3758, 
    3759, 
    3760, 
    3761, 
    3762, 
    3763, 
    3764, 
    3765, 
    3766, 
    3767, 
    3768, 
    3769, 
    3770, 
    3771, 
    3772, 
    3773, 
    3774, 
    3775, 
    3776, 
    3777, 
    3778, 
    3779, 
    3780, 
    3781, 
    3782, 
    3783, 
    3784, 
    3785, 
    3786, 
    3787, 
    3788, 
    3789, 
    3790, 
    3791, 
    3792, 
    3793, 
    3794, 
    3795, 
    3796, 
    3797, 
    3798, 
    3799, 
    3800, 
    3801, 
    3802, 
    3803, 
    3804, 
    3805, 
    3806, 
    3807, 
    3808, 
    3809, 
    3810, 
    3811, 
    3812, 
    3813, 
    3814, 
    3815, 
    3816, 
    3817, 
    3818, 
    3819, 
    3820, 
    3821, 
    3822, 
    3823, 
    3824, 
    3825, 
    3826, 
    3827, 
    3828, 
    3829, 
    3830, 
    3831, 
    3832, 
    3833, 
    3834, 
    3835, 
    3836, 
    3837, 
    3838, 
    3839, 
    3840, 
    3841, 
    3842, 
    3843, 
    3844, 
    3845, 
    3846, 
    3847, 
    3848, 
    3849, 
    3850, 
    3851, 
    3852, 
    3853, 
    3854, 
    3855, 
    3856, 
    3857, 
    3858, 
    3859, 
    3860, 
    3861, 
    3862, 
    3863, 
    3864, 
    3865, 
    3866, 
    3867, 
    3868, 
    3869, 
    3870, 
    3871, 
    3872, 
    3873, 
    3874, 
    3875, 
    3876, 
    3877, 
    3878, 
    3879, 
    3880, 
    3881, 
    3882, 
    3883, 
    3884, 
    3885, 
    3886, 
    3887, 
    3888, 
    3889, 
    3890, 
    3891, 
    3892, 
    3893, 
    3894, 
    3895, 
    3896, 
    3897, 
    3898, 
    3899, 
    3900, 
    3901, 
    3902, 
    3903, 
    3904, 
    3905, 
    3906, 
    3907, 
    3908, 
    3909, 
    3910, 
    3911, 
    3912, 
    3913, 
    3914, 
    3915, 
    3916, 
    3917, 
    3918, 
    3919, 
    3920, 
    3921, 
    3922, 
    3923, 
    3924, 
    3925, 
    3926, 
    3927, 
    3928, 
    3929, 
    3930, 
    3931, 
    3932, 
    3933, 
    3934, 
    3935, 
    3936, 
    3937, 
    3938, 
    3939, 
    3940, 
    3941, 
    3942, 
    3943, 
    3944, 
    3945, 
    3946, 
    3947, 
    3948, 
    3949, 
    3950, 
    3951, 
    3952, 
    3953, 
    3954, 
    3955, 
    3956, 
    3957, 
    3958, 
    3959, 
    3960, 
    3961, 
    3962, 
    3963, 
    3964, 
    3965, 
    3966, 
    3967, 
    3968, 
    3969, 
    3970, 
    3971, 
    3972, 
    3973, 
    3974, 
    3975, 
    3976, 
    3977, 
    3978, 
    3979, 
    3980, 
    3981, 
    3982, 
    3983, 
    3984, 
    3985, 
    3986, 
    3987, 
    3988, 
    3989, 
    3990, 
    3991, 
    3992, 
    3993, 
    3994, 
    3995, 
    3996, 
    3997, 
    3998, 
    3999, 
    4000, 
    4001, 
    4002, 
    4003, 
    4004, 
    4005, 
    4006, 
    4007, 
    4008, 
    4009, 
    4010, 
    4011, 
    4012, 
    4013, 
    4014, 
    4015, 
    4016, 
    4017, 
    4018, 
    4019, 
    4020, 
    4021, 
    4022, 
    4023, 
    4024, 
    4025, 
    4026, 
    4027, 
    4028, 
    4029, 
    4030, 
    4031, 
    4032, 
    4033, 
    4034, 
    4035, 
    4036, 
    4037, 
    4038, 
    4039, 
    4040, 
    4041, 
    4042, 
    4043, 
    4044, 
    4045, 
    4046, 
    4047, 
    4048, 
    4049, 
    4050, 
    4051, 
    4052, 
    4053, 
    4054, 
    4055, 
    4056, 
    4057, 
    4058, 
    4059, 
    4060, 
    4061, 
    4062, 
    4063, 
    4064, 
    4065, 
    4066, 
    4067, 
    4068, 
    4069, 
    4070, 
    4071, 
    4072, 
    4073, 
    4074, 
    4075, 
    4076, 
    4077, 
    4078, 
    4079, 
    4080, 
    4081, 
    4082, 
    4083, 
    4084, 
    4085, 
    4086, 
    4087, 
    4088, 
    4089, 
    4090, 
    4091, 
    4092, 
    4093, 
    4094, 
    4095, 
    4096, 
    4097, 
    4098, 
    4099, 
    4100, 
    4101, 
    4102, 
    4103, 
    4104, 
    4105, 
    4106, 
    4107, 
    4108, 
    4109, 
    4110, 
    4111, 
    4112, 
    4113, 
    4114, 
    4115, 
    4116, 
    4117, 
    4118, 
    4119, 
    4120, 
    4121, 
    4122, 
    4123, 
    4124, 
    4125, 
    4126, 
    4127, 
    4128, 
    4129, 
    4130, 
    4131, 
    4132, 
    4133, 
    4134, 
    4135, 
    4136, 
    4137, 
    4138, 
    4139, 
    4140, 
    4141, 
    4142, 
    4143, 
    4144, 
    4145, 
    4146, 
    4147, 
    4148, 
    4149, 
    4150, 
    4151, 
    4152, 
    4153, 
    4154, 
    4155, 
    4156, 
    4157, 
    4158, 
    4159, 
    4160, 
    4161, 
    4162, 
    4163, 
    4164, 
    4165, 
    4166, 
    4167, 
    4168, 
    4169, 
    4170, 
    4171, 
    4172, 
    4173, 
    4174, 
    4175, 
    4176, 
    4177, 
    4178, 
    4179, 
    4180, 
    4181, 
    4182, 
    4183, 
    4184, 
    4185, 
    4186, 
    4187, 
    4188, 
    4189, 
    4190, 
    4191, 
    4192, 
    4193, 
    4194, 
    4195, 
    4196, 
    4197, 
    4198, 
    4199, 
    4200, 
    4201, 
    4202, 
    4203, 
    4204, 
    4205, 
    4206, 
    4207, 
    4208, 
    4209, 
    4210, 
    4211, 
    4212, 
    4213, 
    4214, 
    4215, 
    4216, 
    4217, 
    4218, 
    4219, 
    4220, 
    4221, 
    4222, 
    4223, 
    4224, 
    4225, 
    4226, 
    4227, 
    4228, 
    4229, 
    4230, 
    4231, 
    4232, 
    4233, 
    4234, 
    4235, 
    4236, 
    4237, 
    4238, 
    4239, 
    4240, 
    4241, 
    4242, 
    4243, 
    4244, 
    4245, 
    4246, 
    4247, 
    4248, 
    4249, 
    4250, 
    4251, 
    4252, 
    4253, 
    4254, 
    4255, 
    4256, 
    4257, 
    4258, 
    4259, 
    4260, 
    4261, 
    4262, 
    4263, 
    4264, 
    4265, 
    4266, 
    4267, 
    4268, 
    4269, 
    4270, 
    4271, 
    4272, 
    4273, 
    4274, 
    4275, 
    4276, 
    4277, 
    4278, 
    4279, 
    4280, 
    4281, 
    4282, 
    4283, 
    4284, 
    4285, 
    4286, 
    4287, 
    4288, 
    4289, 
    4290, 
    4291, 
    4292, 
    4293, 
    4294, 
    4295, 
    4296, 
    4297, 
    4298, 
    4299, 
    4300, 
    4301, 
    4302, 
    4303, 
    4304, 
    4305, 
    4306, 
    4307, 
    4308, 
    4309, 
    4310, 
    4311, 
    4312, 
    4313, 
    4314, 
    4315, 
    4316, 
    4317, 
    4318, 
    4319, 
    4320, 
    4321, 
    4322, 
    4323, 
    4324, 
    4325, 
    4326, 
    4327, 
    4328, 
    4329, 
    4330, 
    4331, 
    4332, 
    4333, 
    4334, 
    4335, 
    4336, 
    4337, 
    4338, 
    4339, 
    4340, 
    4341, 
    4342, 
    4343, 
    4344, 
    4345, 
    4346, 
    4347, 
    4348, 
    4349, 
    4350, 
    4351, 
    4352, 
    4353, 
    4354, 
    4355, 
    4356, 
    4357, 
    4358, 
    4359, 
    4360, 
    4361, 
    4362, 
    4363, 
    4364, 
    4365, 
    4366, 
    4367, 
    4368, 
    4369, 
    4370, 
    4371, 
    4372, 
    4373, 
    4374, 
    4375, 
    4376, 
    4377, 
    4378, 
    4379, 
    4380, 
    4381, 
    4382, 
    4383, 
    4384, 
    4385, 
    4386, 
    4387, 
    4388, 
    4389, 
    4390, 
    4391, 
    4392, 
    4393, 
    4394, 
    4395, 
    4396, 
    4397, 
    4398, 
    4399, 
    4400, 
    4401, 
    4402, 
    4403, 
    4404, 
    4405, 
    4406, 
    4407, 
    4408, 
    4409, 
    4410, 
    4411, 
    4412, 
    4413, 
    4414, 
    4415, 
    4416, 
    4417, 
    4418, 
    4419, 
    4420, 
    4421, 
    4422, 
    4423, 
    4424, 
    4425, 
    4426, 
    4427, 
    4428, 
    4429, 
    4430, 
    4431, 
    4432, 
    4433, 
    4434, 
    4435, 
    4436, 
    4437, 
    4438, 
    4439, 
    4440, 
    4441, 
    4442, 
    4443, 
    4444, 
    4445, 
    4446, 
    4447, 
    4448, 
    4449, 
    4450, 
    4451, 
    4452, 
    4453, 
    4454, 
    4455, 
    4456, 
    4457, 
    4458, 
    4459, 
    4460, 
    4461, 
    4462, 
    4463, 
    4464, 
    4465, 
    4466, 
    4467, 
    4468, 
    4469, 
    4470, 
    4471, 
    4472, 
    4473, 
    4474, 
    4475, 
    4476, 
    4477, 
    4478, 
    4479, 
    4480, 
    4481, 
    4482, 
    4483, 
    4484, 
    4485, 
    4486, 
    4487, 
    4488, 
    4489, 
    4490, 
    4491, 
    4492, 
    4493, 
    4494, 
    4495, 
    4496, 
    4497, 
    4498, 
    4499, 
    4500, 
    4501, 
    4502, 
    4503, 
    4504, 
    4505, 
    4506, 
    4507, 
    4508, 
    4509, 
    4510, 
    4511, 
    4512, 
    4513, 
    4514, 
    4515, 
    4516, 
    4517, 
    4518, 
    4519, 
    4520, 
    4521, 
    4522, 
    4523, 
    4524, 
    4525, 
    4526, 
    4527, 
    4528, 
    4529, 
    4530, 
    4531, 
    4532, 
    4533, 
    4534, 
    4535, 
    4536, 
    4537, 
    4538, 
    4539, 
    4540, 
    4541, 
    4542, 
    4543, 
    4544, 
    4545, 
    4546, 
    4547, 
    4548, 
    4549, 
    4550, 
    4551, 
    4552, 
    4553, 
    4554, 
    4555, 
    4556, 
    4557, 
    4558, 
    4559, 
    4560, 
    4561, 
    4562, 
    4563, 
    4564, 
    4565, 
    4566, 
    4567, 
    4568, 
    4569, 
    4570, 
    4571, 
    4572, 
    4573, 
    4574, 
    4575, 
    4576, 
    4577, 
    4578, 
    4579, 
    4580, 
    4581, 
    4582, 
    4583, 
    4584, 
    4585, 
    4586, 
    4587, 
    4588, 
    4589, 
    4590, 
    4591, 
    4592, 
    4593, 
    4594, 
    4595, 
    4596, 
    4597, 
    4598, 
    4599, 
    4600, 
    4601, 
    4602, 
    4603, 
    4604, 
    4605, 
    4606, 
    4607, 
    4608, 
    4609, 
    4610, 
    4611, 
    4612, 
    4613, 
    4614, 
    4615, 
    4616, 
    4617, 
    4618, 
    4619, 
    4620, 
    4621, 
    4622, 
    4623, 
    4624, 
    4625, 
    4626, 
    4627, 
    4628, 
    4629, 
    4630, 
    4631, 
    4632, 
    4633, 
    4634, 
    4635, 
    4636, 
    4637, 
    4638, 
    4639, 
    4640, 
    4641, 
    4642, 
    4643, 
    4644, 
    4645, 
    4646, 
    4647, 
    4648, 
    4649, 
    4650, 
    4651, 
    4652, 
    4653, 
    4654, 
    4655, 
    4656, 
    4657, 
    4658, 
    4659, 
    4660, 
    4661, 
    4662, 
    4663, 
    4664, 
    4665, 
    4666, 
    4667, 
    4668, 
    4669, 
    4670, 
    4671, 
    4672, 
    4673, 
    4674, 
    4675, 
    4676, 
    4677, 
    4678, 
    4679, 
    4680, 
    4681, 
    4682, 
    4683, 
    4684, 
    4685, 
    4686, 
    4687, 
    4688, 
    4689, 
    4690, 
    4691, 
    4692, 
    4693, 
    4694, 
    4695, 
    4696, 
    4697, 
    4698, 
    4699, 
    4700, 
    4701, 
    4702, 
    4703, 
    4704, 
    4705, 
    4706, 
    4707, 
    4708, 
    4709, 
    4710, 
    4711, 
    4712, 
    4713, 
    4714, 
    4715, 
    4716, 
    4717, 
    4718, 
    4719, 
    4720, 
    4721, 
    4722, 
    4723, 
    4724, 
    4725, 
    4726, 
    4727, 
    4728, 
    4729, 
    4730, 
    4731, 
    4732, 
    4733, 
    4734, 
    4735, 
    4736, 
    4737, 
    4738, 
    4739, 
    4740, 
    4741, 
    4742, 
    4743, 
    4744, 
    4745, 
    4746, 
    4747, 
    4748, 
    4749, 
    4750, 
    4751, 
    4752, 
    4753, 
    4754, 
    4755, 
    4756, 
    4757, 
    4758, 
    4759, 
    4760, 
    4761, 
    4762, 
    4763, 
    4764, 
    4765, 
    4766, 
    4767, 
    4768, 
    4769, 
    4770, 
    4771, 
    4772, 
    4773, 
    4774, 
    4775, 
    4776, 
    4777, 
    4778, 
    4779, 
    4780, 
    4781, 
    4782, 
    4783, 
    4784, 
    4785, 
    4786, 
    4787, 
    4788, 
    4789, 
    4790, 
    4791, 
    4792, 
    4793, 
    4794, 
    4795, 
    4796, 
    4797, 
    4798, 
    4799, 
    4800, 
    4801, 
    4802, 
    4803, 
    4804, 
    4805, 
    4806, 
    4807, 
    4808, 
    4809, 
    4810, 
    4811, 
    4812, 
    4813, 
    4814, 
    4815, 
    4816, 
    4817, 
    4818, 
    4819, 
    4820, 
    4821, 
    4822, 
    4823, 
    4824, 
    4825, 
    4826, 
    4827, 
    4828, 
    4829, 
    4830, 
    4831, 
    4832, 
    4833, 
    4834, 
    4835, 
    4836, 
    4837, 
    4838, 
    4839, 
    4840, 
    4841, 
    4842, 
    4843, 
    4844, 
    4845, 
    4846, 
    4847, 
    4848, 
    4849, 
    4850, 
    4851, 
    4852, 
    4853, 
    4854, 
    4855, 
    4856, 
    4857, 
    4858, 
    4859, 
    4860, 
    4861, 
    4862, 
    4863, 
    4864, 
    4865, 
    4866, 
    4867, 
    4868, 
    4869, 
    4870, 
    4871, 
    4872, 
    4873, 
    4874, 
    4875, 
    4876, 
    4877, 
    4878, 
    4879, 
    4880, 
    4881, 
    4882, 
    4883, 
    4884, 
    4885, 
    4886, 
    4887, 
    4888, 
    4889, 
    4890, 
    4891, 
    4892, 
    4893, 
    4894, 
    4895, 
    4896, 
    4897, 
    4898, 
    4899, 
    4900, 
    4901, 
    4902, 
    4903, 
    4904, 
    4905, 
    4906, 
    4907, 
    4908, 
    4909, 
    4910, 
    4911, 
    4912, 
    4913, 
    4914, 
    4915, 
    4916, 
    4917, 
    4918, 
    4919, 
    4920, 
    4921, 
    4922, 
    4923, 
    4924, 
    4925, 
    4926, 
    4927, 
    4928, 
    4929, 
    4930, 
    4931, 
    4932, 
    4933, 
    4934, 
    4935, 
    4936, 
    4937, 
    4938, 
    4939, 
    4940, 
    4941, 
    4942, 
    4943, 
    4944, 
    4945, 
    4946, 
    4947, 
    4948, 
    4949, 
    4950, 
    4951, 
    4952, 
    4953, 
    4954, 
    4955, 
    4956, 
    4957, 
    4958, 
    4959, 
    4960, 
    4961, 
    4962, 
    4963, 
    4964, 
    4965, 
    4966, 
    4967, 
    4968, 
    4969, 
    4970, 
    4971, 
    4972, 
    4973, 
    4974, 
    4975, 
    4976, 
    4977, 
    4978, 
    4979, 
    4980, 
    4981, 
    4982, 
    4983, 
    4984, 
    4985, 
    4986, 
    4987, 
    4988, 
    4989, 
    4990, 
    4991, 
    4992, 
    4993, 
    4994, 
    4995, 
    4996, 
    4997, 
    4998, 
    4999, 
    5000, 
    5001, 
    5002, 
    5003, 
    5004, 
    5005, 
    5006, 
    5007, 
    5008, 
    5009, 
    5010, 
    5011, 
    5012, 
    5013, 
    5014, 
    5015, 
    5016, 
    5017, 
    5018, 
    5019, 
    5020, 
    5021, 
    5022, 
    5023, 
    5024, 
    5025, 
    5026, 
    5027, 
    5028, 
    5029, 
    5030, 
    5031, 
    5032, 
    5033, 
    5034, 
    5035, 
    5036, 
    5037, 
    5038, 
    5039, 
    5040, 
    5041, 
    5042, 
    5043, 
    5044, 
    5045, 
    5046, 
    5047, 
    5048, 
    5049, 
    5050, 
    5051, 
    5052, 
    5053, 
    5054, 
    5055, 
    5056, 
    5057, 
    5058, 
    5059, 
    5060, 
    5061, 
    5062, 
    5063, 
    5064, 
    5065, 
    5066, 
    5067, 
    5068, 
    5069, 
    5070, 
    5071, 
    5072, 
    5073, 
    5074, 
    5075, 
    5076, 
    5077, 
    5078, 
    5079, 
    5080, 
    5081, 
    5082, 
    5083, 
    5084, 
    5085, 
    5086, 
    5087, 
    5088, 
    5089, 
    5090, 
    5091, 
    5092, 
    5093, 
    5094, 
    5095, 
    5096, 
    5097, 
    5098, 
    5099, 
    5100, 
    5101, 
    5102, 
    5103, 
    5104, 
    5105, 
    5106, 
    5107, 
    5108, 
    5109, 
    5110, 
    5111, 
    5112, 
    5113, 
    5114, 
    5115, 
    5116, 
    5117, 
    5118, 
    5119, 
    5120, 
    5121, 
    5122, 
    5123, 
    5124, 
    5125, 
    5126, 
    5127, 
    5128, 
    5129, 
    5130, 
    5131, 
    5132, 
    5133, 
    5134, 
    5135, 
    5136, 
    5137, 
    5138, 
    5139, 
    5140, 
    5141, 
    5142, 
    5143, 
    5144, 
    5145, 
    5146, 
    5147, 
    5148, 
    5149, 
    5150, 
    5151, 
    5152, 
    5153, 
    5154, 
    5155, 
    5156, 
    5157, 
    5158, 
    5159, 
    5160, 
    5161, 
    5162, 
    5163, 
    5164, 
    5165, 
    5166, 
    5167, 
    5168, 
    5169, 
    5170, 
    5171, 
    5172, 
    5173, 
    5174, 
    5175, 
    5176, 
    5177, 
    5178, 
    5179, 
    5180, 
    5181, 
    5182, 
    5183, 
    5184, 
    5185, 
    5186, 
    5187, 
    5188, 
    5189, 
    5190, 
    5191, 
    5192, 
    5193, 
    5194, 
    5195, 
    5196, 
    5197, 
    5198, 
    5199, 
    5200, 
    5201, 
    5202, 
    5203, 
    5204, 
    5205, 
    5206, 
    5207, 
    5208, 
    5209, 
    5210, 
    5211, 
    5212, 
    5213, 
    5214, 
    5215, 
    5216, 
    5217, 
    5218, 
    5219, 
    5220, 
    5221, 
    5222, 
    5223, 
    5224, 
    5225, 
    5226, 
    5227, 
    5228, 
    5229, 
    5230, 
    5231, 
    5232, 
    5233, 
    5234, 
    5235, 
    5236, 
    5237, 
    5238, 
    5239, 
    5240, 
    5241, 
    5242, 
    5243, 
    5244, 
    5245, 
    5246, 
    5247, 
    5248, 
    5249, 
    5250, 
    5251, 
    5252, 
    5253, 
    5254, 
    5255, 
    5256, 
    5257, 
    5258, 
    5259, 
    5260, 
    5261, 
    5262, 
    5263, 
    5264, 
    5265, 
    5266, 
    5267, 
    5268, 
    5269, 
    5270, 
    5271, 
    5272, 
    5273, 
    5274, 
    5275, 
    5276, 
    5277, 
    5278, 
    5279, 
    5280, 
    5281, 
    5282, 
    5283, 
    5284, 
    5285, 
    5286, 
    5287, 
    5288, 
    5289, 
    5290, 
    5291, 
    5292, 
    5293, 
    5294, 
    5295, 
    5296, 
    5297, 
    5298, 
    5299, 
    5300, 
    5301, 
    5302, 
    5303, 
    5304, 
    5305, 
    5306, 
    5307, 
    5308, 
    5309, 
    5310, 
    5311, 
    5312, 
    5313, 
    5314, 
    5315, 
    5316, 
    5317, 
    5318, 
    5319, 
    5320, 
    5321, 
    5322, 
    5323, 
    5324, 
    5325, 
    5326, 
    5327, 
    5328, 
    5329, 
    5330, 
    5331, 
    5332, 
    5333, 
    5334, 
    5335, 
    5336, 
    5337, 
    5338, 
    5339, 
    5340, 
    5341, 
    5342, 
    5343, 
    5344, 
    5345, 
    5346, 
    5347, 
    5348, 
    5349, 
    5350, 
    5351, 
    5352, 
    5353, 
    5354, 
    5355, 
    5356, 
    5357, 
    5358, 
    5359, 
    5360, 
    5361, 
    5362, 
    5363, 
    5364, 
    5365, 
    5366, 
    5367, 
    5368, 
    5369, 
    5370, 
    5371, 
    5372, 
    5373, 
    5374, 
    5375, 
    5376, 
    5377, 
    5378, 
    5379, 
    5380, 
    5381, 
    5382, 
    5383, 
    5384, 
    5385, 
    5386, 
    5387, 
    5388, 
    5389, 
    5390, 
    5391, 
    5392, 
    5393, 
    5394, 
    5395, 
    5396, 
    5397, 
    5398, 
    5399, 
    5400, 
    5401, 
    5402, 
    5403, 
    5404, 
    5405, 
    5406, 
    5407, 
    5408, 
    5409, 
    5410, 
    5411, 
    5412, 
    5413, 
    5414, 
    5415, 
    5416, 
    5417, 
    5418, 
    5419, 
    5420, 
    5421, 
    5422, 
    5423, 
    5424, 
    5425, 
    5426, 
    5427, 
    5428, 
    5429, 
    5430, 
    5431, 
    5432, 
    5433, 
    5434, 
    5435, 
    5436, 
    5437, 
    5438, 
    5439, 
    5440, 
    5441, 
    5442, 
    5443, 
    5444, 
    5445, 
    5446, 
    5447, 
    5448, 
    5449, 
    5450, 
    5451, 
    5452, 
    5453, 
    5454, 
    5455, 
    5456, 
    5457, 
    5458, 
    5459, 
    5460, 
    5461, 
    5462, 
    5463, 
    5464, 
    5465, 
    5466, 
    5467, 
    5468, 
    5469, 
    5470, 
    5471, 
    5472, 
    5473, 
    5474, 
    5475, 
    5476, 
    5477, 
    5478, 
    5479, 
    5480, 
    5481, 
    5482, 
    5483, 
    5484, 
    5485, 
    5486, 
    5487, 
    5488, 
    5489, 
    5490, 
    5491, 
    5492, 
    5493, 
    5494, 
    5495, 
    5496, 
    5497, 
    5498, 
    5499, 
    5500, 
    5501, 
    5502, 
    5503, 
    5504, 
    5505, 
    5506, 
    5507, 
    5508, 
    5509, 
    5510, 
    5511, 
    5512, 
    5513, 
    5514, 
    5515, 
    5516, 
    5517, 
    5518, 
    5519, 
    5520, 
    5521, 
    5522, 
    5523, 
    5524, 
    5525, 
    5526, 
    5527, 
    5528, 
    5529, 
    5530, 
    5531, 
    5532, 
    5533, 
    5534, 
    5535, 
    5536, 
    5537, 
    5538, 
    5539, 
    5540, 
    5541, 
    5542, 
    5543, 
    5544, 
    5545, 
    5546, 
    5547, 
    5548, 
    5549, 
    5550, 
    5551, 
    5552, 
    5553, 
    5554, 
    5555, 
    5556, 
    5557, 
    5558, 
    5559, 
    5560, 
    5561, 
    5562, 
    5563, 
    5564, 
    5565, 
    5566, 
    5567, 
    5568, 
    5569, 
    5570, 
    5571, 
    5572, 
    5573, 
    5574, 
    5575, 
    5576, 
    5577, 
    5578, 
    5579, 
    5580, 
    5581, 
    5582, 
    5583, 
    5584, 
    5585, 
    5586, 
    5587, 
    5588, 
    5589, 
    5590, 
    5591, 
    5592, 
    5593, 
    5594, 
    5595, 
    5596, 
    5597, 
    5598, 
    5599, 
    5600, 
    5601, 
    5602, 
    5603, 
    5604, 
    5605, 
    5606, 
    5607, 
    5608, 
    5609, 
    5610, 
    5611, 
    5612, 
    5613, 
    5614, 
    5615, 
    5616, 
    5617, 
    5618, 
    5619, 
    5620, 
    5621, 
    5622, 
    5623, 
    5624, 
    5625, 
    5626, 
    5627, 
    5628, 
    5629, 
    5630, 
    5631, 
    5632, 
    5633, 
    5634, 
    5635, 
    5636, 
    5637, 
    5638, 
    5639, 
    5640, 
    5641, 
    5642, 
    5643, 
    5644, 
    5645, 
    5646, 
    5647, 
    5648, 
    5649, 
    5650, 
    5651, 
    5652, 
    5653, 
    5654, 
    5655, 
    5656, 
    5657, 
    5658, 
    5659, 
    5660, 
    5661, 
    5662, 
    5663, 
    5664, 
    5665, 
    5666, 
    5667, 
    5668, 
    5669, 
    5670, 
    5671, 
    5672, 
    5673, 
    5674, 
    5675, 
    5676, 
    5677, 
    5678, 
    5679, 
    5680, 
    5681, 
    5682, 
    5683, 
    5684, 
    5685, 
    5686, 
    5687, 
    5688, 
    5689, 
    5690, 
    5691, 
    5692, 
    5693, 
    5694, 
    5695, 
    5696, 
    5697, 
    5698, 
    5699, 
    5700, 
    5701, 
    5702, 
    5703, 
    5704, 
    5705, 
    5706, 
    5707, 
    5708, 
    5709, 
    5710, 
    5711, 
    5712, 
    5713, 
    5714, 
    5715, 
    5716, 
    5717, 
    5718, 
    5719, 
    5720, 
    5721, 
    5722, 
    5723, 
    5724, 
    5725, 
    5726, 
    5727, 
    5728, 
    5729, 
    5730, 
    5731, 
    5732, 
    5733, 
    5734, 
    5735, 
    5736, 
    5737, 
    5738, 
    5739, 
    5740, 
    5741, 
    5742, 
    5743, 
    5744, 
    5745, 
    5746, 
    5747, 
    5748, 
    5749, 
    5750, 
    5751, 
    5752, 
    5753, 
    5754, 
    5755, 
    5756, 
    5757, 
    5758, 
    5759, 
    5760, 
    5761, 
    5762, 
    5763, 
    5764, 
    5765, 
    5766, 
    5767, 
    5768, 
    5769, 
    5770, 
    5771, 
    5772, 
    5773, 
    5774, 
    5775, 
    5776, 
    5777, 
    5778, 
    5779, 
    5780, 
    5781, 
    5782, 
    5783, 
    5784, 
    5785, 
    5786, 
    5787, 
    5788, 
    5789, 
    5790, 
    5791, 
    5792, 
    5793, 
    5794, 
    5795, 
    5796, 
    5797, 
    5798, 
    5799, 
    5800, 
    5801, 
    5802, 
    5803, 
    5804, 
    5805, 
    5806, 
    5807, 
    5808, 
    5809, 
    5810, 
    5811, 
    5812, 
    5813, 
    5814, 
    5815, 
    5816, 
    5817, 
    5818, 
    5819, 
    5820, 
    5821, 
    5822, 
    5823, 
    5824, 
    5825, 
    5826, 
    5827, 
    5828, 
    5829, 
    5830, 
    5831, 
    5832, 
    5833, 
    5834, 
    5835, 
    5836, 
    5837, 
    5838, 
    5839, 
    5840, 
    5841, 
    5842, 
    5843, 
    5844, 
    5845, 
    5846, 
    5847, 
    5848, 
    5849, 
    5850, 
    5851, 
    5852, 
    5853, 
    5854, 
    5855, 
    5856, 
    5857, 
    5858, 
    5859, 
    5860, 
    5861, 
    5862, 
    5863, 
    5864, 
    5865, 
    5866, 
    5867, 
    5868, 
    5869, 
    5870, 
    5871, 
    5872, 
    5873, 
    5874, 
    5875, 
    5876, 
    5877, 
    5878, 
    5879, 
    5880, 
    5881, 
    5882, 
    5883, 
    5884, 
    5885, 
    5886, 
    5887, 
    5888, 
    5889, 
    5890, 
    5891, 
    5892, 
    5893, 
    5894, 
    5895, 
    5896, 
    5897, 
    5898, 
    5899, 
    5900, 
    5901, 
    5902, 
    5903, 
    5904, 
    5905, 
    5906, 
    5907, 
    5908, 
    5909, 
    5910, 
    5911, 
    5912, 
    5913, 
    5914, 
    5915, 
    5916, 
    5917, 
    5918, 
    5919, 
    5920, 
    5921, 
    5922, 
    5923, 
    5924, 
    5925, 
    5926, 
    5927, 
    5928, 
    5929, 
    5930, 
    5931, 
    5932, 
    5933, 
    5934, 
    5935, 
    5936, 
    5937, 
    5938, 
    5939, 
    5940, 
    5941, 
    5942, 
    5943, 
    5944, 
    5945, 
    5946, 
    5947, 
    5948, 
    5949, 
    5950, 
    5951, 
    5952, 
    5953, 
    5954, 
    5955, 
    5956, 
    5957, 
    5958, 
    5959, 
    5960, 
    5961, 
    5962, 
    5963, 
    5964, 
    5965, 
    5966, 
    5967, 
    5968, 
    5969, 
    5970, 
    5971, 
    5972, 
    5973, 
    5974, 
    5975, 
    5976, 
    5977, 
    5978, 
    5979, 
    5980, 
    5981, 
    5982, 
    5983, 
    5984, 
    5985, 
    5986, 
    5987, 
    5988, 
    5989, 
    5990, 
    5991, 
    5992, 
    5993, 
    5994, 
    5995, 
    5996, 
    5997, 
    5998, 
    5999, 
    6000, 
    6001, 
    6002, 
    6003, 
    6004, 
    6005, 
    6006, 
    6007, 
    6008, 
    6009, 
    6010, 
    6011, 
    6012, 
    6013, 
    6014, 
    6015, 
    6016, 
    6017, 
    6018, 
    6019, 
    6020, 
    6021, 
    6022, 
    6023, 
    6024, 
    6025, 
    6026, 
    6027, 
    6028, 
    6029, 
    6030, 
    6031, 
    6032, 
    6033, 
    6034, 
    6035, 
    6036, 
    6037, 
    6038, 
    6039, 
    6040, 
    6041, 
    6042, 
    6043, 
    6044, 
    6045, 
    6046, 
    6047, 
    6048, 
    6049, 
    6050, 
    6051, 
    6052, 
    6053, 
    6054, 
    6055, 
    6056, 
    6057, 
    6058, 
    6059, 
    6060, 
    6061, 
    6062, 
    6063, 
    6064, 
    6065, 
    6066, 
    6067, 
    6068, 
    6069, 
    6070, 
    6071, 
    6072, 
    6073, 
    6074, 
    6075, 
    6076, 
    6077, 
    6078, 
    6079, 
    6080, 
    6081, 
    6082, 
    6083, 
    6084, 
    6085, 
    6086, 
    6087, 
    6088, 
    6089, 
    6090, 
    6091, 
    6092, 
    6093, 
    6094, 
    6095, 
    6096, 
    6097, 
    6098, 
    6099, 
    6100, 
    6101, 
    6102, 
    6103, 
    6104, 
    6105, 
    6106, 
    6107, 
    6108, 
    6109, 
    6110, 
    6111, 
    6112, 
    6113, 
    6114, 
    6115, 
    6116, 
    6117, 
    6118, 
    6119, 
    6120, 
    6121, 
    6122, 
    6123, 
    6124, 
    6125, 
    6126, 
    6127, 
    6128, 
    6129, 
    6130, 
    6131, 
    6132, 
    6133, 
    6134, 
    6135, 
    6136, 
    6137, 
    6138, 
    6139, 
    6140, 
    6141, 
    6142, 
    6143, 
    6144, 
    6145, 
    6146, 
    6147, 
    6148, 
    6149, 
    6150, 
    6151, 
    6152, 
    6153, 
    6154, 
    6155, 
    6156, 
    6157, 
    6158, 
    6159, 
    6160, 
    6161, 
    6162, 
    6163, 
    6164, 
    6165, 
    6166, 
    6167, 
    6168, 
    6169, 
    6170, 
    6171, 
    6172, 
    6173, 
    6174, 
    6175, 
    6176, 
    6177, 
    6178, 
    6179, 
    6180, 
    6181, 
    6182, 
    6183, 
    6184, 
    6185, 
    6186, 
    6187, 
    6188, 
    6189, 
    6190, 
    6191, 
    6192, 
    6193, 
    6194, 
    6195, 
    6196, 
    6197, 
    6198, 
    6199, 
    6200, 
    6201, 
    6202, 
    6203, 
    6204, 
    6205, 
    6206, 
    6207, 
    6208, 
    6209, 
    6210, 
    6211, 
    6212, 
    6213, 
    6214, 
    6215, 
    6216, 
    6217, 
    6218, 
    6219, 
    6220, 
    6221, 
    6222, 
    6223, 
    6224, 
    6225, 
    6226, 
    6227, 
    6228, 
    6229, 
    6230, 
    6231, 
    6232, 
    6233, 
    6234, 
    6235, 
    6236, 
    6237, 
    6238, 
    6239, 
    6240, 
    6241, 
    6242, 
    6243, 
    6244, 
    6245, 
    6246, 
    6247, 
    6248, 
    6249, 
    6250, 
    6251, 
    6252, 
    6253, 
    6254, 
    6255, 
    6256, 
    6257, 
    6258, 
    6259, 
    6260, 
    6261, 
    6262, 
    6263, 
    6264, 
    6265, 
    6266, 
    6267, 
    6268, 
    6269, 
    6270, 
    6271, 
    6272, 
    6273, 
    6274, 
    6275, 
    6276, 
    6277, 
    6278, 
    6279, 
    6280, 
    6281, 
    6282, 
    6283, 
    6284, 
    6285, 
    6286, 
    6287, 
    6288, 
    6289, 
    6290, 
    6291, 
    6292, 
    6293, 
    6294, 
    6295, 
    6296, 
    6297, 
    6298, 
    6299, 
    6300, 
    6301, 
    6302, 
    6303, 
    6304, 
    6305, 
    6306, 
    6307, 
    6308, 
    6309, 
    6310, 
    6311, 
    6312, 
    6313, 
    6314, 
    6315, 
    6316, 
    6317, 
    6318, 
    6319, 
    6320, 
    6321, 
    6322, 
    6323, 
    6324, 
    6325, 
    6326, 
    6327, 
    6328, 
    6329, 
    6330, 
    6331, 
    6332, 
    6333, 
    6334, 
    6335, 
    6336, 
    6337, 
    6338, 
    6339, 
    6340, 
    6341, 
    6342, 
    6343, 
    6344, 
    6345, 
    6346, 
    6347, 
    6348, 
    6349, 
    6350, 
    6351, 
    6352, 
    6353, 
    6354, 
    6355, 
    6356, 
    6357, 
    6358, 
    6359, 
    6360, 
    6361, 
    6362, 
    6363, 
    6364, 
    6365, 
    6366, 
    6367, 
    6368, 
    6369, 
    6370, 
    6371, 
    6372, 
    6373, 
    6374, 
    6375, 
    6376, 
    6377, 
    6378, 
    6379, 
    6380, 
    6381, 
    6382, 
    6383, 
    6384, 
    6385, 
    6386, 
    6387, 
    6388, 
    6389, 
    6390, 
    6391, 
    6392, 
    6393, 
    6394, 
    6395, 
    6396, 
    6397, 
    6398, 
    6399, 
    6400, 
    6401, 
    6402, 
    6403, 
    6404, 
    6405, 
    6406, 
    6407, 
    6408, 
    6409, 
    6410, 
    6411, 
    6412, 
    6413, 
    6414, 
    6415, 
    6416, 
    6417, 
    6418, 
    6419, 
    6420, 
    6421, 
    6422, 
    6423, 
    6424, 
    6425, 
    6426, 
    6427, 
    6428, 
    6429, 
    6430, 
    6431, 
    6432, 
    6433, 
    6434, 
    6435, 
    6436, 
    6437, 
    6438, 
    6439, 
    6440, 
    6441, 
    6442, 
    6443, 
    6444, 
    6445, 
    6446, 
    6447, 
    6448, 
    6449, 
    6450, 
    6451, 
    6452, 
    6453, 
    6454, 
    6455, 
    6456, 
    6457, 
    6458, 
    6459, 
    6460, 
    6461, 
    6462, 
    6463, 
    6464, 
    6465, 
    6466, 
    6467, 
    6468, 
    6469, 
    6470, 
    6471, 
    6472, 
    6473, 
    6474, 
    6475, 
    6476, 
    6477, 
    6478, 
    6479, 
    6480, 
    6481, 
    6482, 
    6483, 
    6484, 
    6485, 
    6486, 
    6487, 
    6488, 
    6489, 
    6490, 
    6491, 
    6492, 
    6493, 
    6494, 
    6495, 
    6496, 
    6497, 
    6498, 
    6499, 
    6500, 
    6501, 
    6502, 
    6503, 
    6504, 
    6505, 
    6506, 
    6507, 
    6508, 
    6509, 
    6510, 
    6511, 
    6512, 
    6513, 
    6514, 
    6515, 
    6516, 
    6517, 
    6518, 
    6519, 
    6520, 
    6521, 
    6522, 
    6523, 
    6524, 
    6525, 
    6526, 
    6527, 
    6528, 
    6529, 
    6530, 
    6531, 
    6532, 
    6533, 
    6534, 
    6535, 
    6536, 
    6537, 
    6538, 
    6539, 
    6540, 
    6541, 
    6542, 
    6543, 
    6544, 
    6545, 
    6546, 
    6547, 
    6548, 
    6549, 
    6550, 
    6551, 
    6552, 
    6553, 
    6554, 
    6555, 
    6556, 
    6557, 
    6558, 
    6559, 
    6560, 
    6561, 
    6562, 
    6563, 
    6564, 
    6565, 
    6566, 
    6567, 
    6568, 
    6569, 
    6570, 
    6571, 
    6572, 
    6573, 
    6574, 
    6575, 
    6576, 
    6577, 
    6578, 
    6579, 
    6580, 
    6581, 
    6582, 
    6583, 
    6584, 
    6585, 
    6586, 
    6587, 
    6588, 
    6589, 
    6590, 
    6591, 
    6592, 
    6593, 
    6594, 
    6595, 
    6596, 
    6597, 
    6598, 
    6599, 
    6600, 
    6601, 
    6602, 
    6603, 
    6604, 
    6605, 
    6606, 
    6607, 
    6608, 
    6609, 
    6610, 
    6611, 
    6612, 
    6613, 
    6614, 
    6615, 
    6616, 
    6617, 
    6618, 
    6619, 
    6620, 
    6621, 
    6622, 
    6623, 
    6624, 
    6625, 
    6626, 
    6627, 
    6628, 
    6629, 
    6630, 
    6631, 
    6632, 
    6633, 
    6634, 
    6635, 
    6636, 
    6637, 
    6638, 
    6639, 
    6640, 
    6641, 
    6642, 
    6643, 
    6644, 
    6645, 
    6646, 
    6647, 
    6648, 
    6649, 
    6650, 
    6651, 
    6652, 
    6653, 
    6654, 
    6655, 
    6656, 
    6657, 
    6658, 
    6659, 
    6660, 
    6661, 
    6662, 
    6663, 
    6664, 
    6665, 
    6666, 
    6667, 
    6668, 
    6669, 
    6670, 
    6671, 
    6672, 
    6673, 
    6674, 
    6675, 
    6676, 
    6677, 
    6678, 
    6679, 
    6680, 
    6681, 
    6682, 
    6683, 
    6684, 
    6685, 
    6686, 
    6687, 
    6688, 
    6689, 
    6690, 
    6691, 
    6692, 
    6693, 
    6694, 
    6695, 
    6696, 
    6697, 
    6698, 
    6699, 
    6700, 
    6701, 
    6702, 
    6703, 
    6704, 
    6705, 
    6706, 
    6707, 
    6708, 
    6709, 
    6710, 
    6711, 
    6712, 
    6713, 
    6714, 
    6715, 
    6716, 
    6717, 
    6718, 
    6719, 
    6720, 
    6721, 
    6722, 
    6723, 
    6724, 
    6725, 
    6726, 
    6727, 
    6728, 
    6729, 
    6730, 
    6731, 
    6732, 
    6733, 
    6734, 
    6735, 
    6736, 
    6737, 
    6738, 
    6739, 
    6740, 
    6741, 
    6742, 
    6743, 
    6744, 
    6745, 
    6746, 
    6747, 
    6748, 
    6749, 
    6750, 
    6751, 
    6752, 
    6753, 
    6754, 
    6755, 
    6756, 
    6757, 
    6758, 
    6759, 
    6760, 
    6761, 
    6762, 
    6763, 
    6764, 
    6765, 
    6766, 
    6767, 
    6768, 
    6769, 
    6770, 
    6771, 
    6772, 
    6773, 
    6774, 
    6775, 
    6776, 
    6777, 
    6778, 
    6779, 
    6780, 
    6781, 
    6782, 
    6783, 
    6784, 
    6785, 
    6786, 
    6787, 
    6788, 
    6789, 
    6790, 
    6791, 
    6792, 
    6793, 
    6794, 
    6795, 
    6796, 
    6797, 
    6798, 
    6799, 
    6800, 
    6801, 
    6802, 
    6803, 
    6804, 
    6805, 
    6806, 
    6807, 
    6808, 
    6809, 
    6810, 
    6811, 
    6812, 
    6813, 
    6814, 
    6815, 
    6816, 
    6817, 
    6818, 
    6819, 
    6820, 
    6821, 
    6822, 
    6823, 
    6824, 
    6825, 
    6826, 
    6827, 
    6828, 
    6829, 
    6830, 
    6831, 
    6832, 
    6833, 
    6834, 
    6835, 
    6836, 
    6837, 
    6838, 
    6839, 
    6840, 
    6841, 
    6842, 
    6843, 
    6844, 
    6845, 
    6846, 
    6847, 
    6848, 
    6849, 
    6850, 
    6851, 
    6852, 
    6853, 
    6854, 
    6855, 
    6856, 
    6857, 
    6858, 
    6859, 
    6860, 
    6861, 
    6862, 
    6863, 
    6864, 
    6865, 
    6866, 
    6867, 
    6868, 
    6869, 
    6870, 
    6871, 
    6872, 
    6873, 
    6874, 
    6875, 
    6876, 
    6877, 
    6878, 
    6879, 
    6880, 
    6881, 
    6882, 
    6883, 
    6884, 
    6885, 
    6886, 
    6887, 
    6888, 
    6889, 
    6890, 
    6891, 
    6892, 
    6893, 
    6894, 
    6895, 
    6896, 
    6897, 
    6898, 
    6899, 
    6900, 
    6901, 
    6902, 
    6903, 
    6904, 
    6905, 
    6906, 
    6907, 
    6908, 
    6909, 
    6910, 
    6911, 
    6912, 
    6913, 
    6914, 
    6915, 
    6916, 
    6917, 
    6918, 
    6919, 
    6920, 
    6921, 
    6922, 
    6923, 
    6924, 
    6925, 
    6926, 
    6927, 
    6928, 
    6929, 
    6930, 
    6931, 
    6932, 
    6933, 
    6934, 
    6935, 
    6936, 
    6937, 
    6938, 
    6939, 
    6940, 
    6941, 
    6942, 
    6943, 
    6944, 
    6945, 
    6946, 
    6947, 
    6948, 
    6949, 
    6950, 
    6951, 
    6952, 
    6953, 
    6954, 
    6955, 
    6956, 
    6957, 
    6958, 
    6959, 
    6960, 
    6961, 
    6962, 
    6963, 
    6964, 
    6965, 
    6966, 
    6967, 
    6968, 
    6969, 
    6970, 
    6971, 
    6972, 
    6973, 
    6974, 
    6975, 
    6976, 
    6977, 
    6978, 
    6979, 
    6980, 
    6981, 
    6982, 
    6983, 
    6984, 
    6985, 
    6986, 
    6987, 
    6988, 
    6989, 
    6990, 
    6991, 
    6992, 
    6993, 
    6994, 
    6995, 
    6996, 
    6997, 
    6998, 
    6999, 
    7000, 
    7001, 
    7002, 
    7003, 
    7004, 
    7005, 
    7006, 
    7007, 
    7008, 
    7009, 
    7010, 
    7011, 
    7012, 
    7013, 
    7014, 
    7015, 
    7016, 
    7017, 
    7018, 
    7019, 
    7020, 
    7021, 
    7022, 
    7023, 
    7024, 
    7025, 
    7026, 
    7027, 
    7028, 
    7029, 
    7030, 
    7031, 
    7032, 
    7033, 
    7034, 
    7035, 
    7036, 
    7037, 
    7038, 
    7039, 
    7040, 
    7041, 
    7042, 
    7043, 
    7044, 
    7045, 
    7046, 
    7047, 
    7048, 
    7049, 
    7050, 
    7051, 
    7052, 
    7053, 
    7054, 
    7055, 
    7056, 
    7057, 
    7058, 
    7059, 
    7060, 
    7061, 
    7062, 
    7063, 
    7064, 
    7065, 
    7066, 
    7067, 
    7068, 
    7069, 
    7070, 
    7071, 
    7072, 
    7073, 
    7074, 
    7075, 
    7076, 
    7077, 
    7078, 
    7079, 
    7080, 
    7081, 
    7082, 
    7083, 
    7084, 
    7085, 
    7086, 
    7087, 
    7088, 
    7089, 
    7090, 
    7091, 
    7092, 
    7093, 
    7094, 
    7095, 
    7096, 
    7097, 
    7098, 
    7099, 
    7100, 
    7101, 
    7102, 
    7103, 
    7104, 
    7105, 
    7106, 
    7107, 
    7108, 
    7109, 
    7110, 
    7111, 
    7112, 
    7113, 
    7114, 
    7115, 
    7116, 
    7117, 
    7118, 
    7119, 
    7120, 
    7121, 
    7122, 
    7123, 
    7124, 
    7125, 
    7126, 
    7127, 
    7128, 
    7129, 
    7130, 
    7131, 
    7132, 
    7133, 
    7134, 
    7135, 
    7136, 
    7137, 
    7138, 
    7139, 
    7140, 
    7141, 
    7142, 
    7143, 
    7144, 
    7145, 
    7146, 
    7147, 
    7148, 
    7149, 
    7150, 
    7151, 
    7152, 
    7153, 
    7154, 
    7155, 
    7156, 
    7157, 
    7158, 
    7159, 
    7160, 
    7161, 
    7162, 
    7163, 
    7164, 
    7165, 
    7166, 
    7167, 
    7168, 
    7169, 
    7170, 
    7171, 
    7172, 
    7173, 
    7174, 
    7175, 
    7176, 
    7177, 
    7178, 
    7179, 
    7180, 
    7181, 
    7182, 
    7183, 
    7184, 
    7185, 
    7186, 
    7187, 
    7188, 
    7189, 
    7190, 
    7191, 
    7192, 
    7193, 
    7194, 
    7195, 
    7196, 
    7197, 
    7198, 
    7199, 
    7200, 
    7201, 
    7202, 
    7203, 
    7204, 
    7205, 
    7206, 
    7207, 
    7208, 
    7209, 
    7210, 
    7211, 
    7212, 
    7213, 
    7214, 
    7215, 
    7216, 
    7217, 
    7218, 
    7219, 
    7220, 
    7221, 
    7222, 
    7223, 
    7224, 
    7225, 
    7226, 
    7227, 
    7228, 
    7229, 
    7230, 
    7231, 
    7232, 
    7233, 
    7234, 
    7235, 
    7236, 
    7237, 
    7238, 
    7239, 
    7240, 
    7241, 
    7242, 
    7243, 
    7244, 
    7245, 
    7246, 
    7247, 
    7248, 
    7249, 
    7250, 
    7251, 
    7252, 
    7253, 
    7254, 
    7255, 
    7256, 
    7257, 
    7258, 
    7259, 
    7260, 
    7261, 
    7262, 
    7263, 
    7264, 
    7265, 
    7266, 
    7267, 
    7268, 
    7269, 
    7270, 
    7271, 
    7272, 
    7273, 
    7274, 
    7275, 
    7276, 
    7277, 
    7278, 
    7279, 
    7280, 
    7281, 
    7282, 
    7283, 
    7284, 
    7285, 
    7286, 
    7287, 
    7288, 
    7289, 
    7290, 
    7291, 
    7292, 
    7293, 
    7294, 
    7295, 
    7296, 
    7297, 
    7298, 
    7299, 
    7300, 
    7301, 
    7302, 
    7303, 
    7304, 
    7305, 
    7306, 
    7307, 
    7308, 
    7309, 
    7310, 
    7311, 
    7312, 
    7313, 
    7314, 
    7315, 
    7316, 
    7317, 
    7318, 
    7319, 
    7320, 
    7321, 
    7322, 
    7323, 
    7324, 
    7325, 
    7326, 
    7327, 
    7328, 
    7329, 
    7330, 
    7331, 
    7332, 
    7333, 
    7334, 
    7335, 
    7336, 
    7337, 
    7338, 
    7339, 
    7340, 
    7341, 
    7342, 
    7343, 
    7344, 
    7345, 
    7346, 
    7347, 
    7348, 
    7349, 
    7350, 
    7351, 
    7352, 
    7353, 
    7354, 
    7355, 
    7356, 
    7357, 
    7358, 
    7359, 
    7360, 
    7361, 
    7362, 
    7363, 
    7364, 
    7365, 
    7366, 
    7367, 
    7368, 
    7369, 
    7370, 
    7371, 
    7372, 
    7373, 
    7374, 
    7375, 
    7376, 
    7377, 
    7378, 
    7379, 
    7380, 
    7381, 
    7382, 
    7383, 
    7384, 
    7385, 
    7386, 
    7387, 
    7388, 
    7389, 
    7390, 
    7391, 
    7392, 
    7393, 
    7394, 
    7395, 
    7396, 
    7397, 
    7398, 
    7399, 
    7400, 
    7401, 
    7402, 
    7403, 
    7404, 
    7405, 
    7406, 
    7407, 
    7408, 
    7409, 
    7410, 
    7411, 
    7412, 
    7413, 
    7414, 
    7415, 
    7416, 
    7417, 
    7418, 
    7419, 
    7420, 
    7421, 
    7422, 
    7423, 
    7424, 
    7425, 
    7426, 
    7427, 
    7428, 
    7429, 
    7430, 
    7431, 
    7432, 
    7433, 
    7434, 
    7435, 
    7436, 
    7437, 
    7438, 
    7439, 
    7440, 
    7441, 
    7442, 
    7443, 
    7444, 
    7445, 
    7446, 
    7447, 
    7448, 
    7449, 
    7450, 
    7451, 
    7452, 
    7453, 
    7454, 
    7455, 
    7456, 
    7457, 
    7458, 
    7459, 
    7460, 
    7461, 
    7462, 
    7463, 
    7464, 
    7465, 
    7466, 
    7467, 
    7468, 
    7469, 
    7470, 
    7471, 
    7472, 
    7473, 
    7474, 
    7475, 
    7476, 
    7477, 
    7478, 
    7479, 
    7480, 
    7481, 
    7482, 
    7483, 
    7484, 
    7485, 
    7486, 
    7487, 
    7488, 
    7489, 
    7490, 
    7491, 
    7492, 
    7493, 
    7494, 
    7495, 
    7496, 
    7497, 
    7498, 
    7499, 
    7500, 
    7501, 
    7502, 
    7503, 
    7504, 
    7505, 
    7506, 
    7507, 
    7508, 
    7509, 
    7510, 
    7511, 
    7512, 
    7513, 
    7514, 
    7515, 
    7516, 
    7517, 
    7518, 
    7519, 
    7520, 
    7521, 
    7522, 
    7523, 
    7524, 
    7525, 
    7526, 
    7527, 
    7528, 
    7529, 
    7530, 
    7531, 
    7532, 
    7533, 
    7534, 
    7535, 
    7536, 
    7537, 
    7538, 
    7539, 
    7540, 
    7541, 
    7542, 
    7543, 
    7544, 
    7545, 
    7546, 
    7547, 
    7548, 
    7549, 
    7550, 
    7551, 
    7552, 
    7553, 
    7554, 
    7555, 
    7556, 
    7557, 
    7558, 
    7559, 
    7560, 
    7561, 
    7562, 
    7563, 
    7564, 
    7565, 
    7566, 
    7567, 
    7568, 
    7569, 
    7570, 
    7571, 
    7572, 
    7573, 
    7574, 
    7575, 
    7576, 
    7577, 
    7578, 
    7579, 
    7580, 
    7581, 
    7582, 
    7583, 
    7584, 
    7585, 
    7586, 
    7587, 
    7588, 
    7589, 
    7590, 
    7591, 
    7592, 
    7593, 
    7594, 
    7595, 
    7596, 
    7597, 
    7598, 
    7599, 
    7600, 
    7601, 
    7602, 
    7603, 
    7604, 
    7605, 
    7606, 
    7607, 
    7608, 
    7609, 
    7610, 
    7611, 
    7612, 
    7613, 
    7614, 
    7615, 
    7616, 
    7617, 
    7618, 
    7619, 
    7620, 
    7621, 
    7622, 
    7623, 
    7624, 
    7625, 
    7626, 
    7627, 
    7628, 
    7629, 
    7630, 
    7631, 
    7632, 
    7633, 
    7634, 
    7635, 
    7636, 
    7637, 
    7638, 
    7639, 
    7640, 
    7641, 
    7642, 
    7643, 
    7644, 
    7645, 
    7646, 
    7647, 
    7648, 
    7649, 
    7650, 
    7651, 
    7652, 
    7653, 
    7654, 
    7655, 
    7656, 
    7657, 
    7658, 
    7659, 
    7660, 
    7661, 
    7662, 
    7663, 
    7664, 
    7665, 
    7666, 
    7667, 
    7668, 
    7669, 
    7670, 
    7671, 
    7672, 
    7673, 
    7674, 
    7675, 
    7676, 
    7677, 
    7678, 
    7679, 
    7680, 
    7681, 
    7682, 
    7683, 
    7684, 
    7685, 
    7686, 
    7687, 
    7688, 
    7689, 
    7690, 
    7691, 
    7692, 
    7693, 
    7694, 
    7695, 
    7696, 
    7697, 
    7698, 
    7699, 
    7700, 
    7701, 
    7702, 
    7703, 
    7704, 
    7705, 
    7706, 
    7707, 
    7708, 
    7709, 
    7710, 
    7711, 
    7712, 
    7713, 
    7714, 
    7715, 
    7716, 
    7717, 
    7718, 
    7719, 
    7720, 
    7721, 
    7722, 
    7723, 
    7724, 
    7725, 
    7726, 
    7727, 
    7728, 
    7729, 
    7730, 
    7731, 
    7732, 
    7733, 
    7734, 
    7735, 
    7736, 
    7737, 
    7738, 
    7739, 
    7740, 
    7741, 
    7742, 
    7743, 
    7744, 
    7745, 
    7746, 
    7747, 
    7748, 
    7749, 
    7750, 
    7751, 
    7752, 
    7753, 
    7754, 
    7755, 
    7756, 
    7757, 
    7758, 
    7759, 
    7760, 
    7761, 
    7762, 
    7763, 
    7764, 
    7765, 
    7766, 
    7767, 
    7768, 
    7769, 
    7770, 
    7771, 
    7772, 
    7773, 
    7774, 
    7775, 
    7776, 
    7777, 
    7778, 
    7779, 
    7780, 
    7781, 
    7782, 
    7783, 
    7784, 
    7785, 
    7786, 
    7787, 
    7788, 
    7789, 
    7790, 
    7791, 
    7792, 
    7793, 
    7794, 
    7795, 
    7796, 
    7797, 
    7798, 
    7799, 
    7800, 
    7801, 
    7802, 
    7803, 
    7804, 
    7805, 
    7806, 
    7807, 
    7808, 
    7809, 
    7810, 
    7811, 
    7812, 
    7813, 
    7814, 
    7815, 
    7816, 
    7817, 
    7818, 
    7819, 
    7820, 
    7821, 
    7822, 
    7823, 
    7824, 
    7825, 
    7826, 
    7827, 
    7828, 
    7829, 
    7830, 
    7831, 
    7832, 
    7833, 
    7834, 
    7835, 
    7836, 
    7837, 
    7838, 
    7839, 
    7840, 
    7841, 
    7842, 
    7843, 
    7844, 
    7845, 
    7846, 
    7847, 
    7848, 
    7849, 
    7850, 
    7851, 
    7852, 
    7853, 
    7854, 
    7855, 
    7856, 
    7857, 
    7858, 
    7859, 
    7860, 
    7861, 
    7862, 
    7863, 
    7864, 
    7865, 
    7866, 
    7867, 
    7868, 
    7869, 
    7870, 
    7871, 
    7872, 
    7873, 
    7874, 
    7875, 
    7876, 
    7877, 
    7878, 
    7879, 
    7880, 
    7881, 
    7882, 
    7883, 
    7884, 
    7885, 
    7886, 
    7887, 
    7888, 
    7889, 
    7890, 
    7891, 
    7892, 
    7893, 
    7894, 
    7895, 
    7896, 
    7897, 
    7898, 
    7899, 
    7900, 
    7901, 
    7902, 
    7903, 
    7904, 
    7905, 
    7906, 
    7907, 
    7908, 
    7909, 
    7910, 
    7911, 
    7912, 
    7913, 
    7914, 
    7915, 
    7916, 
    7917, 
    7918, 
    7919, 
    7920, 
    7921, 
    7922, 
    7923, 
    7924, 
    7925, 
    7926, 
    7927, 
    7928, 
    7929, 
    7930, 
    7931, 
    7932, 
    7933, 
    7934, 
    7935, 
    7936, 
    7937, 
    7938, 
    7939, 
    7940, 
    7941, 
    7942, 
    7943, 
    7944, 
    7945, 
    7946, 
    7947, 
    7948, 
    7949, 
    7950, 
    7951, 
    7952, 
    7953, 
    7954, 
    7955, 
    7956, 
    7957, 
    7958, 
    7959, 
    7960, 
    7961, 
    7962, 
    7963, 
    7964, 
    7965, 
    7966, 
    7967, 
    7968, 
    7969, 
    7970, 
    7971, 
    7972, 
    7973, 
    7974, 
    7975, 
    7976, 
    7977, 
    7978, 
    7979, 
    7980, 
    7981, 
    7982, 
    7983, 
    7984, 
    7985, 
    7986, 
    7987, 
    7988, 
    7989, 
    7990, 
    7991, 
    7992, 
    7993, 
    7994, 
    7995, 
    7996, 
    7997, 
    7998, 
    7999, 
    8000, 
    8001, 
    8002, 
    8003, 
    8004, 
    8005, 
    8006, 
    8007, 
    8008, 
    8009, 
    8010, 
    8011, 
    8012, 
    8013, 
    8014, 
    8015, 
    8016, 
    8017, 
    8018, 
    8019, 
    8020, 
    8021, 
    8022, 
    8023, 
    8024, 
    8025, 
    8026, 
    8027, 
    8028, 
    8029, 
    8030, 
    8031, 
    8032, 
    8033, 
    8034, 
    8035, 
    8036, 
    8037, 
    8038, 
    8039, 
    8040, 
    8041, 
    8042, 
    8043, 
    8044, 
    8045, 
    8046, 
    8047, 
    8048, 
    8049, 
    8050, 
    8051, 
    8052, 
    8053, 
    8054, 
    8055, 
    8056, 
    8057, 
    8058, 
    8059, 
    8060, 
    8061, 
    8062, 
    8063, 
    8064, 
    8065, 
    8066, 
    8067, 
    8068, 
    8069, 
    8070, 
    8071, 
    8072, 
    8073, 
    8074, 
    8075, 
    8076, 
    8077, 
    8078, 
    8079, 
    8080, 
    8081, 
    8082, 
    8083, 
    8084, 
    8085, 
    8086, 
    8087, 
    8088, 
    8089, 
    8090, 
    8091, 
    8092, 
    8093, 
    8094, 
    8095, 
    8096, 
    8097, 
    8098, 
    8099, 
    8100, 
    8101, 
    8102, 
    8103, 
    8104, 
    8105, 
    8106, 
    8107, 
    8108, 
    8109, 
    8110, 
    8111, 
    8112, 
    8113, 
    8114, 
    8115, 
    8116, 
    8117, 
    8118, 
    8119, 
    8120, 
    8121, 
    8122, 
    8123, 
    8124, 
    8125, 
    8126, 
    8127, 
    8128, 
    8129, 
    8130, 
    8131, 
    8132, 
    8133, 
    8134, 
    8135, 
    8136, 
    8137, 
    8138, 
    8139, 
    8140, 
    8141, 
    8142, 
    8143, 
    8144, 
    8145, 
    8146, 
    8147, 
    8148, 
    8149, 
    8150, 
    8151, 
    8152, 
    8153, 
    8154, 
    8155, 
    8156, 
    8157, 
    8158, 
    8159, 
    8160, 
    8161, 
    8162, 
    8163, 
    8164, 
    8165, 
    8166, 
    8167, 
    8168, 
    8169, 
    8170, 
    8171, 
    8172, 
    8173, 
    8174, 
    8175, 
    8176, 
    8177, 
    8178, 
    8179, 
    8180, 
    8181, 
    8182, 
    8183, 
    8184, 
    8185, 
    8186, 
    8187, 
    8188, 
    8189, 
    8190, 
    8191, 
    8192, 
    8193, 
    8194, 
    8195, 
    8196, 
    8197, 
    8198, 
    8199, 
    8200, 
    8201, 
    8202, 
    8203, 
    8204, 
    8205, 
    8206, 
    8207, 
    8208, 
    8209, 
    8210, 
    8211, 
    8212, 
    8213, 
    8214, 
    8215, 
    8216, 
    8217, 
    8218, 
    8219, 
    8220, 
    8221, 
    8222, 
    8223, 
    8224, 
    8225, 
    8226, 
    8227, 
    8228, 
    8229, 
    8230, 
    8231, 
    8232, 
    8233, 
    8234, 
    8235, 
    8236, 
    8237, 
    8238, 
    8239, 
    8240, 
    8241, 
    8242, 
    8243, 
    8244, 
    8245, 
    8246, 
    8247, 
    8248, 
    8249, 
    8250, 
    8251, 
    8252, 
    8253, 
    8254, 
    8255, 
    8256, 
    8257, 
    8258, 
    8259, 
    8260, 
    8261, 
    8262, 
    8263, 
    8264, 
    8265, 
    8266, 
    8267, 
    8268, 
    8269, 
    8270, 
    8271, 
    8272, 
    8273, 
    8274, 
    8275, 
    8276, 
    8277, 
    8278, 
    8279, 
    8280, 
    8281, 
    8282, 
    8283, 
    8284, 
    8285, 
    8286, 
    8287, 
    8288, 
    8289, 
    8290, 
    8291, 
    8292, 
    8293, 
    8294, 
    8295, 
    8296, 
    8297, 
    8298, 
    8299, 
    8300, 
    8301, 
    8302, 
    8303, 
    8304, 
    8305, 
    8306, 
    8307, 
    8308, 
    8309, 
    8310, 
    8311, 
    8312, 
    8313, 
    8314, 
    8315, 
    8316, 
    8317, 
    8318, 
    8319, 
    8320, 
    8321, 
    8322, 
    8323, 
    8324, 
    8325, 
    8326, 
    8327, 
    8328, 
    8329, 
    8330, 
    8331, 
    8332, 
    8333, 
    8334, 
    8335, 
    8336, 
    8337, 
    8338, 
    8339, 
    8340, 
    8341, 
    8342, 
    8343, 
    8344, 
    8345, 
    8346, 
    8347, 
    8348, 
    8349, 
    8350, 
    8351, 
    8352, 
    8353, 
    8354, 
    8355, 
    8356, 
    8357, 
    8358, 
    8359, 
    8360, 
    8361, 
    8362, 
    8363, 
    8364, 
    8365, 
    8366, 
    8367, 
    8368, 
    8369, 
    8370, 
    8371, 
    8372, 
    8373, 
    8374, 
    8375, 
    8376, 
    8377, 
    8378, 
    8379, 
    8380, 
    8381, 
    8382, 
    8383, 
    8384, 
    8385, 
    8386, 
    8387, 
    8388, 
    8389, 
    8390, 
    8391, 
    8392, 
    8393, 
    8394, 
    8395, 
    8396, 
    8397, 
    8398, 
    8399, 
    8400, 
    8401, 
    8402, 
    8403, 
    8404, 
    8405, 
    8406, 
    8407, 
    8408, 
    8409, 
    8410, 
    8411, 
    8412, 
    8413, 
    8414, 
    8415, 
    8416, 
    8417, 
    8418, 
    8419, 
    8420, 
    8421, 
    8422, 
    8423, 
    8424, 
    8425, 
    8426, 
    8427, 
    8428, 
    8429, 
    8430, 
    8431, 
    8432, 
    8433, 
    8434, 
    8435, 
    8436, 
    8437, 
    8438, 
    8439, 
    8440, 
    8441, 
    8442, 
    8443, 
    8444, 
    8445, 
    8446, 
    8447, 
    8448, 
    8449, 
    8450, 
    8451, 
    8452, 
    8453, 
    8454, 
    8455, 
    8456, 
    8457, 
    8458, 
    8459, 
    8460, 
    8461, 
    8462, 
    8463, 
    8464, 
    8465, 
    8466, 
    8467, 
    8468, 
    8469, 
    8470, 
    8471, 
    8472, 
    8473, 
    8474, 
    8475, 
    8476, 
    8477, 
    8478, 
    8479, 
    8480, 
    8481, 
    8482, 
    8483, 
    8484, 
    8485, 
    8486, 
    8487, 
    8488, 
    8489, 
    8490, 
    8491, 
    8492, 
    8493, 
    8494, 
    8495, 
    8496, 
    8497, 
    8498, 
    8499, 
    8500, 
    8501, 
    8502, 
    8503, 
    8504, 
    8505, 
    8506, 
    8507, 
    8508, 
    8509, 
    8510, 
    8511, 
    8512, 
    8513, 
    8514, 
    8515, 
    8516, 
    8517, 
    8518, 
    8519, 
    8520, 
    8521, 
    8522, 
    8523, 
    8524, 
    8525, 
    8526, 
    8527, 
    8528, 
    8529, 
    8530, 
    8531, 
    8532, 
    8533, 
    8534, 
    8535, 
    8536, 
    8537, 
    8538, 
    8539, 
    8540, 
    8541, 
    8542, 
    8543, 
    8544, 
    8545, 
    8546, 
    8547, 
    8548, 
    8549, 
    8550, 
    8551, 
    8552, 
    8553, 
    8554, 
    8555, 
    8556, 
    8557, 
    8558, 
    8559, 
    8560, 
    8561, 
    8562, 
    8563, 
    8564, 
    8565, 
    8566, 
    8567, 
    8568, 
    8569, 
    8570, 
    8571, 
    8572, 
    8573, 
    8574, 
    8575, 
    8576, 
    8577, 
    8578, 
    8579, 
    8580, 
    8581, 
    8582, 
    8583, 
    8584, 
    8585, 
    8586, 
    8587, 
    8588, 
    8589, 
    8590, 
    8591, 
    8592, 
    8593, 
    8594, 
    8595, 
    8596, 
    8597, 
    8598, 
    8599, 
    8600, 
    8601, 
    8602, 
    8603, 
    8604, 
    8605, 
    8606, 
    8607, 
    8608, 
    8609, 
    8610, 
    8611, 
    8612, 
    8613, 
    8614, 
    8615, 
    8616, 
    8617, 
    8618, 
    8619, 
    8620, 
    8621, 
    8622, 
    8623, 
    8624, 
    8625, 
    8626, 
    8627, 
    8628, 
    8629, 
    8630, 
    8631, 
    8632, 
    8633, 
    8634, 
    8635, 
    8636, 
    8637, 
    8638, 
    8639, 
    8640, 
    8641, 
    8642, 
    8643, 
    8644, 
    8645, 
    8646, 
    8647, 
    8648, 
    8649, 
    8650, 
    8651, 
    8652, 
    8653, 
    8654, 
    8655, 
    8656, 
    8657, 
    8658, 
    8659, 
    8660, 
    8661, 
    8662, 
    8663, 
    8664, 
    8665, 
    8666, 
    8667, 
    8668, 
    8669, 
    8670, 
    8671, 
    8672, 
    8673, 
    8674, 
    8675, 
    8676, 
    8677, 
    8678, 
    8679, 
    8680, 
    8681, 
    8682, 
    8683, 
    8684, 
    8685, 
    8686, 
    8687, 
    8688, 
    8689, 
    8690, 
    8691, 
    8692, 
    8693, 
    8694, 
    8695, 
    8696, 
    8697, 
    8698, 
    8699, 
    8700, 
    8701, 
    8702, 
    8703, 
    8704, 
    8705, 
    8706, 
    8707, 
    8708, 
    8709, 
    8710, 
    8711, 
    8712, 
    8713, 
    8714, 
    8715, 
    8716, 
    8717, 
    8718, 
    8719, 
    8720, 
    8721, 
    8722, 
    8723, 
    8724, 
    8725, 
    8726, 
    8727, 
    8728, 
    8729, 
    8730, 
    8731, 
    8732, 
    8733, 
    8734, 
    8735, 
    8736, 
    8737, 
    8738, 
    8739, 
    8740, 
    8741, 
    8742, 
    8743, 
    8744, 
    8745, 
    8746, 
    8747, 
    8748, 
    8749, 
    8750, 
    8751, 
    8752, 
    8753, 
    8754, 
    8755, 
    8756, 
    8757, 
    8758, 
    8759, 
    8760, 
    8761, 
    8762, 
    8763, 
    8764, 
    8765, 
    8766, 
    8767, 
    8768, 
    8769, 
    8770, 
    8771, 
    8772, 
    8773, 
    8774, 
    8775, 
    8776, 
    8777, 
    8778, 
    8779, 
    8780, 
    8781, 
    8782, 
    8783, 
    8784, 
    8785, 
    8786, 
    8787, 
    8788, 
    8789, 
    8790, 
    8791, 
    8792, 
    8793, 
    8794, 
    8795, 
    8796, 
    8797, 
    8798, 
    8799, 
    8800, 
    8801, 
    8802, 
    8803, 
    8804, 
    8805, 
    8806, 
    8807, 
    8808, 
    8809, 
    8810, 
    8811, 
    8812, 
    8813, 
    8814, 
    8815, 
    8816, 
    8817, 
    8818, 
    8819, 
    8820, 
    8821, 
    8822, 
    8823, 
    8824, 
    8825, 
    8826, 
    8827, 
    8828, 
    8829, 
    8830, 
    8831, 
    8832, 
    8833, 
    8834, 
    8835, 
    8836, 
    8837, 
    8838, 
    8839, 
    8840, 
    8841, 
    8842, 
    8843, 
    8844, 
    8845, 
    8846, 
    8847, 
    8848, 
    8849, 
    8850, 
    8851, 
    8852, 
    8853, 
    8854, 
    8855, 
    8856, 
    8857, 
    8858, 
    8859, 
    8860, 
    8861, 
    8862, 
    8863, 
    8864, 
    8865, 
    8866, 
    8867, 
    8868, 
    8869, 
    8870, 
    8871, 
    8872, 
    8873, 
    8874, 
    8875, 
    8876, 
    8877, 
    8878, 
    8879, 
    8880, 
    8881, 
    8882, 
    8883, 
    8884, 
    8885, 
    8886, 
    8887, 
    8888, 
    8889, 
    8890, 
    8891, 
    8892, 
    8893, 
    8894, 
    8895, 
    8896, 
    8897, 
    8898, 
    8899, 
    8900, 
    8901, 
    8902, 
    8903, 
    8904, 
    8905, 
    8906, 
    8907, 
    8908, 
    8909, 
    8910, 
    8911, 
    8912, 
    8913, 
    8914, 
    8915, 
    8916, 
    8917, 
    8918, 
    8919, 
    8920, 
    8921, 
    8922, 
    8923, 
    8924, 
    8925, 
    8926, 
    8927, 
    8928, 
    8929, 
    8930, 
    8931, 
    8932, 
    8933, 
    8934, 
    8935, 
    8936, 
    8937, 
    8938, 
    8939, 
    8940, 
    8941, 
    8942, 
    8943, 
    8944, 
    8945, 
    8946, 
    8947, 
    8948, 
    8949, 
    8950, 
    8951, 
    8952, 
    8953, 
    8954, 
    8955, 
    8956, 
    8957, 
    8958, 
    8959, 
    8960, 
    8961, 
    8962, 
    8963, 
    8964, 
    8965, 
    8966, 
    8967, 
    8968, 
    8969, 
    8970, 
    8971, 
    8972, 
    8973, 
    8974, 
    8975, 
    8976, 
    8977, 
    8978, 
    8979, 
    8980, 
    8981, 
    8982, 
    8983, 
    8984, 
    8985, 
    8986, 
    8987, 
    8988, 
    8989, 
    8990, 
    8991, 
    8992, 
    8993, 
    8994, 
    8995, 
    8996, 
    8997, 
    8998, 
    8999, 
    9000, 
    9001, 
    9002, 
    9003, 
    9004, 
    9005, 
    9006, 
    9007, 
    9008, 
    9009, 
    9010, 
    9011, 
    9012, 
    9013, 
    9014, 
    9015, 
    9016, 
    9017, 
    9018, 
    9019, 
    9020, 
    9021, 
    9022, 
    9023, 
    9024, 
    9025, 
    9026, 
    9027, 
    9028, 
    9029, 
    9030, 
    9031, 
    9032, 
    9033, 
    9034, 
    9035, 
    9036, 
    9037, 
    9038, 
    9039, 
    9040, 
    9041, 
    9042, 
    9043, 
    9044, 
    9045, 
    9046, 
    9047, 
    9048, 
    9049, 
    9050, 
    9051, 
    9052, 
    9053, 
    9054, 
    9055, 
    9056, 
    9057, 
    9058, 
    9059, 
    9060, 
    9061, 
    9062, 
    9063, 
    9064, 
    9065, 
    9066, 
    9067, 
    9068, 
    9069, 
    9070, 
    9071, 
    9072, 
    9073, 
    9074, 
    9075, 
    9076, 
    9077, 
    9078, 
    9079, 
    9080, 
    9081, 
    9082, 
    9083, 
    9084, 
    9085, 
    9086, 
    9087, 
    9088, 
    9089, 
    9090, 
    9091, 
    9092, 
    9093, 
    9094, 
    9095, 
    9096, 
    9097, 
    9098, 
    9099, 
    9100, 
    9101, 
    9102, 
    9103, 
    9104, 
    9105, 
    9106, 
    9107, 
    9108, 
    9109, 
    9110, 
    9111, 
    9112, 
    9113, 
    9114, 
    9115, 
    9116, 
    9117, 
    9118, 
    9119, 
    9120, 
    9121, 
    9122, 
    9123, 
    9124, 
    9125, 
    9126, 
    9127, 
    9128, 
    9129, 
    9130, 
    9131, 
    9132, 
    9133, 
    9134, 
    9135, 
    9136, 
    9137, 
    9138, 
    9139, 
    9140, 
    9141, 
    9142, 
    9143, 
    9144, 
    9145, 
    9146, 
    9147, 
    9148, 
    9149, 
    9150, 
    9151, 
    9152, 
    9153, 
    9154, 
    9155, 
    9156, 
    9157, 
    9158, 
    9159, 
    9160, 
    9161, 
    9162, 
    9163, 
    9164, 
    9165, 
    9166, 
    9167, 
    9168, 
    9169, 
    9170, 
    9171, 
    9172, 
    9173, 
    9174, 
    9175, 
    9176, 
    9177, 
    9178, 
    9179, 
    9180, 
    9181, 
    9182, 
    9183, 
    9184, 
    9185, 
    9186, 
    9187, 
    9188, 
    9189, 
    9190, 
    9191, 
    9192, 
    9193, 
    9194, 
    9195, 
    9196, 
    9197, 
    9198, 
    9199, 
    9200, 
    9201, 
    9202, 
    9203, 
    9204, 
    9205, 
    9206, 
    9207, 
    9208, 
    9209, 
    9210, 
    9211, 
    9212, 
    9213, 
    9214, 
    9215, 
    9216, 
    9217, 
    9218, 
    9219, 
    9220, 
    9221, 
    9222, 
    9223, 
    9224, 
    9225, 
    9226, 
    9227, 
    9228, 
    9229, 
    9230, 
    9231, 
    9232, 
    9233, 
    9234, 
    9235, 
    9236, 
    9237, 
    9238, 
    9239, 
    9240, 
    9241, 
    9242, 
    9243, 
    9244, 
    9245, 
    9246, 
    9247, 
    9248, 
    9249, 
    9250, 
    9251, 
    9252, 
    9253, 
    9254, 
    9255, 
    9256, 
    9257, 
    9258, 
    9259, 
    9260, 
    9261, 
    9262, 
    9263, 
    9264, 
    9265, 
    9266, 
    9267, 
    9268, 
    9269, 
    9270, 
    9271, 
    9272, 
    9273, 
    9274, 
    9275, 
    9276, 
    9277, 
    9278, 
    9279, 
    9280, 
    9281, 
    9282, 
    9283, 
    9284, 
    9285, 
    9286, 
    9287, 
    9288, 
    9289, 
    9290, 
    9291, 
    9292, 
    9293, 
    9294, 
    9295, 
    9296, 
    9297, 
    9298, 
    9299, 
    9300, 
    9301, 
    9302, 
    9303, 
    9304, 
    9305, 
    9306, 
    9307, 
    9308, 
    9309, 
    9310, 
    9311, 
    9312, 
    9313, 
    9314, 
    9315, 
    9316, 
    9317, 
    9318, 
    9319, 
    9320, 
    9321, 
    9322, 
    9323, 
    9324, 
    9325, 
    9326, 
    9327, 
    9328, 
    9329, 
    9330, 
    9331, 
    9332, 
    9333, 
    9334, 
    9335, 
    9336, 
    9337, 
    9338, 
    9339, 
    9340, 
    9341, 
    9342, 
    9343, 
    9344, 
    9345, 
    9346, 
    9347, 
    9348, 
    9349, 
    9350, 
    9351, 
    9352, 
    9353, 
    9354, 
    9355, 
    9356, 
    9357, 
    9358, 
    9359, 
    9360, 
    9361, 
    9362, 
    9363, 
    9364, 
    9365, 
    9366, 
    9367, 
    9368, 
    9369, 
    9370, 
    9371, 
    9372, 
    9373, 
    9374, 
    9375, 
    9376, 
    9377, 
    9378, 
    9379, 
    9380, 
    9381, 
    9382, 
    9383, 
    9384, 
    9385, 
    9386, 
    9387, 
    9388, 
    9389, 
    9390, 
    9391, 
    9392, 
    9393, 
    9394, 
    9395, 
    9396, 
    9397, 
    9398, 
    9399, 
    9400, 
    9401, 
    9402, 
    9403, 
    9404, 
    9405, 
    9406, 
    9407, 
    9408, 
    9409, 
    9410, 
    9411, 
    9412, 
    9413, 
    9414, 
    9415, 
    9416, 
    9417, 
    9418, 
    9419, 
    9420, 
    9421, 
    9422, 
    9423, 
    9424, 
    9425, 
    9426, 
    9427, 
    9428, 
    9429, 
    9430, 
    9431, 
    9432, 
    9433, 
    9434, 
    9435, 
    9436, 
    9437, 
    9438, 
    9439, 
    9440, 
    9441, 
    9442, 
    9443, 
    9444, 
    9445, 
    9446, 
    9447, 
    9448, 
    9449, 
    9450, 
    9451, 
    9452, 
    9453, 
    9454, 
    9455, 
    9456, 
    9457, 
    9458, 
    9459, 
    9460, 
    9461, 
    9462, 
    9463, 
    9464, 
    9465, 
    9466, 
    9467, 
    9468, 
    9469, 
    9470, 
    9471, 
    9472, 
    9473, 
    9474, 
    9475, 
    9476, 
    9477, 
    9478, 
    9479, 
    9480, 
    9481, 
    9482, 
    9483, 
    9484, 
    9485, 
    9486, 
    9487, 
    9488, 
    9489, 
    9490, 
    9491, 
    9492, 
    9493, 
    9494, 
    9495, 
    9496, 
    9497, 
    9498, 
    9499, 
    9500, 
    9501, 
    9502, 
    9503, 
    9504, 
    9505, 
    9506, 
    9507, 
    9508, 
    9509, 
    9510, 
    9511, 
    9512, 
    9513, 
    9514, 
    9515, 
    9516, 
    9517, 
    9518, 
    9519, 
    9520, 
    9521, 
    9522, 
    9523, 
    9524, 
    9525, 
    9526, 
    9527, 
    9528, 
    9529, 
    9530, 
    9531, 
    9532, 
    9533, 
    9534, 
    9535, 
    9536, 
    9537, 
    9538, 
    9539, 
    9540, 
    9541, 
    9542, 
    9543, 
    9544, 
    9545, 
    9546, 
    9547, 
    9548, 
    9549, 
    9550, 
    9551, 
    9552, 
    9553, 
    9554, 
    9555, 
    9556, 
    9557, 
    9558, 
    9559, 
    9560, 
    9561, 
    9562, 
    9563, 
    9564, 
    9565, 
    9566, 
    9567, 
    9568, 
    9569, 
    9570, 
    9571, 
    9572, 
    9573, 
    9574, 
    9575, 
    9576, 
    9577, 
    9578, 
    9579, 
    9580, 
    9581, 
    9582, 
    9583, 
    9584, 
    9585, 
    9586, 
    9587, 
    9588, 
    9589, 
    9590, 
    9591, 
    9592, 
    9593, 
    9594, 
    9595, 
    9596, 
    9597, 
    9598, 
    9599, 
    9600, 
    9601, 
    9602, 
    9603, 
    9604, 
    9605, 
    9606, 
    9607, 
    9608, 
    9609, 
    9610, 
    9611, 
    9612, 
    9613, 
    9614, 
    9615, 
    9616, 
    9617, 
    9618, 
    9619, 
    9620, 
    9621, 
    9622, 
    9623, 
    9624, 
    9625, 
    9626, 
    9627, 
    9628, 
    9629, 
    9630, 
    9631, 
    9632, 
    9633, 
    9634, 
    9635, 
    9636, 
    9637, 
    9638, 
    9639, 
    9640, 
    9641, 
    9642, 
    9643, 
    9644, 
    9645, 
    9646, 
    9647, 
    9648, 
    9649, 
    9650, 
    9651, 
    9652, 
    9653, 
    9654, 
    9655, 
    9656, 
    9657, 
    9658, 
    9659, 
    9660, 
    9661, 
    9662, 
    9663, 
    9664, 
    9665, 
    9666, 
    9667, 
    9668, 
    9669, 
    9670, 
    9671, 
    9672, 
    9673, 
    9674, 
    9675, 
    9676, 
    9677, 
    9678, 
    9679, 
    9680, 
    9681, 
    9682, 
    9683, 
    9684, 
    9685, 
    9686, 
    9687, 
    9688, 
    9689, 
    9690, 
    9691, 
    9692, 
    9693, 
    9694, 
    9695, 
    9696, 
    9697, 
    9698, 
    9699, 
    9700, 
    9701, 
    9702, 
    9703, 
    9704, 
    9705, 
    9706, 
    9707, 
    9708, 
    9709, 
    9710, 
    9711, 
    9712, 
    9713, 
    9714, 
    9715, 
    9716, 
    9717, 
    9718, 
    9719, 
    9720, 
    9721, 
    9722, 
    9723, 
    9724, 
    9725, 
    9726, 
    9727, 
    9728, 
    9729, 
    9730, 
    9731, 
    9732, 
    9733, 
    9734, 
    9735, 
    9736, 
    9737, 
    9738, 
    9739, 
    9740, 
    9741, 
    9742, 
    9743, 
    9744, 
    9745, 
    9746, 
    9747, 
    9748, 
    9749, 
    9750, 
    9751, 
    9752, 
    9753, 
    9754, 
    9755, 
    9756, 
    9757, 
    9758, 
    9759, 
    9760, 
    9761, 
    9762, 
    9763, 
    9764, 
    9765, 
    9766, 
    9767, 
    9768, 
    9769, 
    9770, 
    9771, 
    9772, 
    9773, 
    9774, 
    9775, 
    9776, 
    9777, 
    9778, 
    9779, 
    9780, 
    9781, 
    9782, 
    9783, 
    9784, 
    9785, 
    9786, 
    9787, 
    9788, 
    9789, 
    9790, 
    9791, 
    9792, 
    9793, 
    9794, 
    9795, 
    9796, 
    9797, 
    9798, 
    9799, 
    9800, 
    9801, 
    9802, 
    9803, 
    9804, 
    9805, 
    9806, 
    9807, 
    9808, 
    9809, 
    9810, 
    9811, 
    9812, 
    9813, 
    9814, 
    9815, 
    9816, 
    9817, 
    9818, 
    9819, 
    9820, 
    9821, 
    9822, 
    9823, 
    9824, 
    9825, 
    9826, 
    9827, 
    9828, 
    9829, 
    9830, 
    9831, 
    9832, 
    9833, 
    9834, 
    9835, 
    9836, 
    9837, 
    9838, 
    9839, 
    9840, 
    9841, 
    9842, 
    9843, 
    9844, 
    9845, 
    9846, 
    9847, 
    9848, 
    9849, 
    9850, 
    9851, 
    9852, 
    9853, 
    9854, 
    9855, 
    9856, 
    9857, 
    9858, 
    9859, 
    9860, 
    9861, 
    9862, 
    9863, 
    9864, 
    9865, 
    9866, 
    9867, 
    9868, 
    9869, 
    9870, 
    9871, 
    9872, 
    9873, 
    9874, 
    9875, 
    9876, 
    9877, 
    9878, 
    9879, 
    9880, 
    9881, 
    9882, 
    9883, 
    9884, 
    9885, 
    9886, 
    9887, 
    9888, 
    9889, 
    9890, 
    9891, 
    9892, 
    9893, 
    9894, 
    9895, 
    9896, 
    9897, 
    9898, 
    9899, 
    9900, 
    9901, 
    9902, 
    9903, 
    9904, 
    9905, 
    9906, 
    9907, 
    9908, 
    9909, 
    9910, 
    9911, 
    9912, 
    9913, 
    9914, 
    9915, 
    9916, 
    9917, 
    9918, 
    9919, 
    9920, 
    9921, 
    9922, 
    9923, 
    9924, 
    9925, 
    9926, 
    9927, 
    9928, 
    9929, 
    9930, 
    9931, 
    9932, 
    9933, 
    9934, 
    9935, 
    9936, 
    9937, 
    9938, 
    9939, 
    9940, 
    9941, 
    9942, 
    9943, 
    9944, 
    9945, 
    9946, 
    9947, 
    9948, 
    9949, 
    9950, 
    9951, 
    9952, 
    9953, 
    9954, 
    9955, 
    9956, 
    9957, 
    9958, 
    9959, 
    9960, 
    9961, 
    9962, 
    9963, 
    9964, 
    9965, 
    9966, 
    9967, 
    9968, 
    9969, 
    9970, 
    9971, 
    9972, 
    9973, 
    9974, 
    9975, 
    9976, 
    9977, 
    9978, 
    9979, 
    9980, 
    9981, 
    9982, 
    9983, 
    9984, 
    9985, 
    9986, 
    9987, 
    9988, 
    9989, 
    9990, 
    9991, 
    9992, 
    9993, 
    9994, 
    9995, 
    9996, 
    9997, 
    9998, 
    9999, 
    10000, 
    10001, 
    10002, 
    10003, 
    10004, 
    10005, 
    10006, 
    10007, 
    10008, 
    10009, 
    10010, 
    10011, 
    10012, 
    10013, 
    10014, 
    10015, 
    10016, 
    10017, 
    10018, 
    10019, 
    10020, 
    10021, 
    10022, 
    10023, 
    10024, 
    10025, 
    10026, 
    10027, 
    10028, 
    10029, 
    10030, 
    10031, 
    10032, 
    10033, 
    10034, 
    10035, 
    10036, 
    10037, 
    10038, 
    10039, 
    10040, 
    10041, 
    10042, 
    10043, 
    10044, 
    10045, 
    10046, 
    10047, 
    10048, 
    10049, 
    10050, 
    10051, 
    10052, 
    10053, 
    10054, 
    10055, 
    10056, 
    10057, 
    10058, 
    10059, 
    10060, 
    10061, 
    10062, 
    10063, 
    10064, 
    10065, 
    10066, 
    10067, 
    10068, 
    10069, 
    10070, 
    10071, 
    10072, 
    10073, 
    10074, 
    10075, 
    10076, 
    10077, 
    10078, 
    10079, 
    10080, 
    10081, 
    10082, 
    10083, 
    10084, 
    10085, 
    10086, 
    10087, 
    10088, 
    10089, 
    10090, 
    10091, 
    10092, 
    10093, 
    10094, 
    10095, 
    10096, 
    10097, 
    10098, 
    10099, 
    10100, 
    10101, 
    10102, 
    10103, 
    10104, 
    10105, 
    10106, 
    10107, 
    10108, 
    10109, 
    10110, 
    10111, 
    10112, 
    10113, 
    10114, 
    10115, 
    10116, 
    10117, 
    10118, 
    10119, 
    10120, 
    10121, 
    10122, 
    10123, 
    10124, 
    10125, 
    10126, 
    10127, 
    10128, 
    10129, 
    10130, 
    10131, 
    10132, 
    10133, 
    10134, 
    10135, 
    10136, 
    10137, 
    10138, 
    10139, 
    10140, 
    10141, 
    10142, 
    10143, 
    10144, 
    10145, 
    10146, 
    10147, 
    10148, 
    10149, 
    10150, 
    10151, 
    10152, 
    10153, 
    10154, 
    10155, 
    10156, 
    10157, 
    10158, 
    10159, 
    10160, 
    10161, 
    10162, 
    10163, 
    10164, 
    10165, 
    10166, 
    10167, 
    10168, 
    10169, 
    10170, 
    10171, 
    10172, 
    10173, 
    10174, 
    10175, 
    10176, 
    10177, 
    10178, 
    10179, 
    10180, 
    10181, 
    10182, 
    10183, 
    10184, 
    10185, 
    10186, 
    10187, 
    10188, 
    10189, 
    10190, 
    10191, 
    10192, 
    10193, 
    10194, 
    10195, 
    10196, 
    10197, 
    10198, 
    10199, 
    10200, 
    10201, 
    10202, 
    10203, 
    10204, 
    10205, 
    10206, 
    10207, 
    10208, 
    10209, 
    10210, 
    10211, 
    10212, 
    10213, 
    10214, 
    10215, 
    10216, 
    10217, 
    10218, 
    10219, 
    10220, 
    10221, 
    10222, 
    10223, 
    10224, 
    10225, 
    10226, 
    10227, 
    10228, 
    10229, 
    10230, 
    10231, 
    10232, 
    10233, 
    10234, 
    10235, 
    10236, 
    10237, 
    10238, 
    10239, 
    10240, 
    10241, 
    10242, 
    10243, 
    10244, 
    10245, 
    10246, 
    10247, 
    10248, 
    10249, 
    10250, 
    10251, 
    10252, 
    10253, 
    10254, 
    10255, 
    10256, 
    10257, 
    10258, 
    10259, 
    10260, 
    10261, 
    10262, 
    10263, 
    10264, 
    10265, 
    10266, 
    10267, 
    10268, 
    10269, 
    10270, 
    10271, 
    10272, 
    10273, 
    10274, 
    10275, 
    10276, 
    10277, 
    10278, 
    10279, 
    10280, 
    10281, 
    10282, 
    10283, 
    10284, 
    10285, 
    10286, 
    10287, 
    10288, 
    10289, 
    10290, 
    10291, 
    10292, 
    10293, 
    10294, 
    10295, 
    10296, 
    10297, 
    10298, 
    10299, 
    10300, 
    10301, 
    10302, 
    10303, 
    10304, 
    10305, 
    10306, 
    10307, 
    10308, 
    10309, 
    10310, 
    10311, 
    10312, 
    10313, 
    10314, 
    10315, 
    10316, 
    10317, 
    10318, 
    10319, 
    10320, 
    10321, 
    10322, 
    10323, 
    10324, 
    10325, 
    10326, 
    10327, 
    10328, 
    10329, 
    10330, 
    10331, 
    10332, 
    10333, 
    10334, 
    10335, 
    10336, 
    10337, 
    10338, 
    10339, 
    10340, 
    10341, 
    10342, 
    10343, 
    10344, 
    10345, 
    10346, 
    10347, 
    10348, 
    10349, 
    10350, 
    10351, 
    10352, 
    10353, 
    10354, 
    10355, 
    10356, 
    10357, 
    10358, 
    10359, 
    10360, 
    10361, 
    10362, 
    10363, 
    10364, 
    10365, 
    10366, 
    10367, 
    10368, 
    10369, 
    10370, 
    10371, 
    10372, 
    10373, 
    10374, 
    10375, 
    10376, 
    10377, 
    10378, 
    10379, 
    10380, 
    10381, 
    10382, 
    10383, 
    10384, 
    10385, 
    10386, 
    10387, 
    10388, 
    10389, 
    10390, 
    10391, 
    10392, 
    10393, 
    10394, 
    10395, 
    10396, 
    10397, 
    10398, 
    10399, 
    10400, 
    10401, 
    10402, 
    10403, 
    10404, 
    10405, 
    10406, 
    10407, 
    10408, 
    10409, 
    10410, 
    10411, 
    10412, 
    10413, 
    10414, 
    10415, 
    10416, 
    10417, 
    10418, 
    10419, 
    10420, 
    10421, 
    10422, 
    10423, 
    10424, 
    10425, 
    10426, 
    10427, 
    10428, 
    10429, 
    10430, 
    10431, 
    10432, 
    10433, 
    10434, 
    10435, 
    10436, 
    10437, 
    10438, 
    10439, 
    10440, 
    10441, 
    10442, 
    10443, 
    10444, 
    10445, 
    10446, 
    10447, 
    10448, 
    10449, 
    10450, 
    10451, 
    10452, 
    10453, 
    10454, 
    10455, 
    10456, 
    10457, 
    10458, 
    10459, 
    10460, 
    10461, 
    10462, 
    10463, 
    10464, 
    10465, 
    10466, 
    10467, 
    10468, 
    10469, 
    10470, 
    10471, 
    10472, 
    10473, 
    10474, 
    10475, 
    10476, 
    10477, 
    10478, 
    10479, 
    10480, 
    10481, 
    10482, 
    10483, 
    10484, 
    10485, 
    10486, 
    10487, 
    10488, 
    10489, 
    10490, 
    10491, 
    10492, 
    10493, 
    10494, 
    10495, 
    10496, 
    10497, 
    10498, 
    10499, 
    10500, 
    10501, 
    10502, 
    10503, 
    10504, 
    10505, 
    10506, 
    10507, 
    10508, 
    10509, 
    10510, 
    10511, 
    10512, 
    10513, 
    10514, 
    10515, 
    10516, 
    10517, 
    10518, 
    10519, 
    10520, 
    10521, 
    10522, 
    10523, 
    10524, 
    10525, 
    10526, 
    10527, 
    10528, 
    10529, 
    10530, 
    10531, 
    10532, 
    10533, 
    10534, 
    10535, 
    10536, 
    10537, 
    10538, 
    10539, 
    10540, 
    10541, 
    10542, 
    10543, 
    10544, 
    10545, 
    10546, 
    10547, 
    10548, 
    10549, 
    10550, 
    10551, 
    10552, 
    10553, 
    10554, 
    10555, 
    10556, 
    10557, 
    10558, 
    10559, 
    10560, 
    10561, 
    10562, 
    10563, 
    10564, 
    10565, 
    10566, 
    10567, 
    10568, 
    10569, 
    10570, 
    10571, 
    10572, 
    10573, 
    10574, 
    10575, 
    10576, 
    10577, 
    10578, 
    10579, 
    10580, 
    10581, 
    10582, 
    10583, 
    10584, 
    10585, 
    10586, 
    10587, 
    10588, 
    10589, 
    10590, 
    10591, 
    10592, 
    10593, 
    10594, 
    10595, 
    10596, 
    10597, 
    10598, 
    10599, 
    10600, 
    10601, 
    10602, 
    10603, 
    10604, 
    10605, 
    10606, 
    10607, 
    10608, 
    10609, 
    10610, 
    10611, 
    10612, 
    10613, 
    10614, 
    10615, 
    10616, 
    10617, 
    10618, 
    10619, 
    10620, 
    10621, 
    10622, 
    10623, 
    10624, 
    10625, 
    10626, 
    10627, 
    10628, 
    10629, 
    10630, 
    10631, 
    10632, 
    10633, 
    10634, 
    10635, 
    10636, 
    10637, 
    10638, 
    10639, 
    10640, 
    10641, 
    10642, 
    10643, 
    10644, 
    10645, 
    10646, 
    10647, 
    10648, 
    10649, 
    10650, 
    10651, 
    10652, 
    10653, 
    10654, 
    10655, 
    10656, 
    10657, 
    10658, 
    10659, 
    10660, 
    10661, 
    10662, 
    10663, 
    10664, 
    10665, 
    10666, 
    10667, 
    10668, 
    10669, 
    10670, 
    10671, 
    10672, 
    10673, 
    10674, 
    10675, 
    10676, 
    10677, 
    10678, 
    10679, 
    10680, 
    10681, 
    10682, 
    10683, 
    10684, 
    10685, 
    10686, 
    10687, 
    10688, 
    10689, 
    10690, 
    10691, 
    10692, 
    10693, 
    10694, 
    10695, 
    10696, 
    10697, 
    10698, 
    10699, 
    10700, 
    10701, 
    10702, 
    10703, 
    10704, 
    10705, 
    10706, 
    10707, 
    10708, 
    10709, 
    10710, 
    10711, 
    10712, 
    10713, 
    10714, 
    10715, 
    10716, 
    10717, 
    10718, 
    10719, 
    10720, 
    10721, 
    10722, 
    10723, 
    10724, 
    10725, 
    10726, 
    10727, 
    10728, 
    10729, 
    10730, 
    10731, 
    10732, 
    10733, 
    10734, 
    10735, 
    10736, 
    10737, 
    10738, 
    10739, 
    10740, 
    10741, 
    10742, 
    10743, 
    10744, 
    10745, 
    10746, 
    10747, 
    10748, 
    10749, 
    10750, 
    10751, 
    10752, 
    10753, 
    10754, 
    10755, 
    10756, 
    10757, 
    10758, 
    10759, 
    10760, 
    10761, 
    10762, 
    10763, 
    10764, 
    10765, 
    10766, 
    10767, 
    10768, 
    10769, 
    10770, 
    10771, 
    10772, 
    10773, 
    10774, 
    10775, 
    10776, 
    10777, 
    10778, 
    10779, 
    10780, 
    10781, 
    10782, 
    10783, 
    10784, 
    10785, 
    10786, 
    10787, 
    10788, 
    10789, 
    10790, 
    10791, 
    10792, 
    10793, 
    10794, 
    10795, 
    10796, 
    10797, 
    10798, 
    10799, 
    10800, 
    10801, 
    10802, 
    10803, 
    10804, 
    10805, 
    10806, 
    10807, 
    10808, 
    10809, 
    10810, 
    10811, 
    10812, 
    10813, 
    10814, 
    10815, 
    10816, 
    10817, 
    10818, 
    10819, 
    10820, 
    10821, 
    10822, 
    10823, 
    10824, 
    10825, 
    10826, 
    10827, 
    10828, 
    10829, 
    10830, 
    10831, 
    10832, 
    10833, 
    10834, 
    10835, 
    10836, 
    10837, 
    10838, 
    10839, 
    10840, 
    10841, 
    10842, 
    10843, 
    10844, 
    10845, 
    10846, 
    10847, 
    10848, 
    10849, 
    10850, 
    10851, 
    10852, 
    10853, 
    10854, 
    10855, 
    10856, 
    10857, 
    10858, 
    10859, 
    10860, 
    10861, 
    10862, 
    10863, 
    10864, 
    10865, 
    10866, 
    10867, 
    10868, 
    10869, 
    10870, 
    10871, 
    10872, 
    10873, 
    10874, 
    10875, 
    10876, 
    10877, 
    10878, 
    10879, 
    10880, 
    10881, 
    10882, 
    10883, 
    10884, 
    10885, 
    10886, 
    10887, 
    10888, 
    10889, 
    10890, 
    10891, 
    10892, 
    10893, 
    10894, 
    10895, 
    10896, 
    10897, 
    10898, 
    10899, 
    10900, 
    10901, 
    10902, 
    10903, 
    10904, 
    10905, 
    10906, 
    10907, 
    10908, 
    10909, 
    10910, 
    10911, 
    10912, 
    10913, 
    10914, 
    10915, 
    10916, 
    10917, 
    10918, 
    10919, 
    10920, 
    10921, 
    10922, 
    10923, 
    10924, 
    10925, 
    10926, 
    10927, 
    10928, 
    10929, 
    10930, 
    10931, 
    10932, 
    10933, 
    10934, 
    10935, 
    10936, 
    10937, 
    10938, 
    10939, 
    10940, 
    10941, 
    10942, 
    10943, 
    10944, 
    10945, 
    10946, 
    10947, 
    10948, 
    10949, 
    10950, 
    10951, 
    10952, 
    10953, 
    10954, 
    10955, 
    10956, 
    10957, 
    10958, 
    10959, 
    10960, 
    10961, 
    10962, 
    10963, 
    10964, 
    10965, 
    10966, 
    10967, 
    10968, 
    10969, 
    10970, 
    10971, 
    10972, 
    10973, 
    10974, 
    10975, 
    10976, 
    10977, 
    10978, 
    10979, 
    10980, 
    10981, 
    10982, 
    10983, 
    10984, 
    10985, 
    10986, 
    10987, 
    10988, 
    10989, 
    10990, 
    10991, 
    10992, 
    10993, 
    10994, 
    10995, 
    10996, 
    10997, 
    10998, 
    10999, 
    11000, 
    11001, 
    11002, 
    11003, 
    11004, 
    11005, 
    11006, 
    11007, 
    11008, 
    11009, 
    11010, 
    11011, 
    11012, 
    11013, 
    11014, 
    11015, 
    11016, 
    11017, 
    11018, 
    11019, 
    11020, 
    11021, 
    11022, 
    11023, 
    11024, 
    11025, 
    11026, 
    11027, 
    11028, 
    11029, 
    11030, 
    11031, 
    11032, 
    11033, 
    11034, 
    11035, 
    11036, 
    11037, 
    11038, 
    11039, 
    11040, 
    11041, 
    11042, 
    11043, 
    11044, 
    11045, 
    11046, 
    11047, 
    11048, 
    11049, 
    11050, 
    11051, 
    11052, 
    11053, 
    11054, 
    11055, 
    11056, 
    11057, 
    11058, 
    11059, 
    11060, 
    11061, 
    11062, 
    11063, 
    11064, 
    11065, 
    11066, 
    11067, 
    11068, 
    11069, 
    11070, 
    11071, 
    11072, 
    11073, 
    11074, 
    11075, 
    11076, 
    11077, 
    11078, 
    11079, 
    11080, 
    11081, 
    11082, 
    11083, 
    11084, 
    11085, 
    11086, 
    11087, 
    11088, 
    11089, 
    11090, 
    11091, 
    11092, 
    11093, 
    11094, 
    11095, 
    11096, 
    11097, 
    11098, 
    11099, 
    11100, 
    11101, 
    11102, 
    11103, 
    11104, 
    11105, 
    11106, 
    11107, 
    11108, 
    11109, 
    11110, 
    11111, 
    11112, 
    11113, 
    11114, 
    11115, 
    11116, 
    11117, 
    11118, 
    11119, 
    11120, 
    11121, 
    11122, 
    11123, 
    11124, 
    11125, 
    11126, 
    11127, 
    11128, 
    11129, 
    11130, 
    11131, 
    11132, 
    11133, 
    11134, 
    11135, 
    11136, 
    11137, 
    11138, 
    11139, 
    11140, 
    11141, 
    11142, 
    11143, 
    11144, 
    11145, 
    11146, 
    11147, 
    11148, 
    11149, 
    11150, 
    11151, 
    11152, 
    11153, 
    11154, 
    11155, 
    11156, 
    11157, 
    11158, 
    11159, 
    11160, 
    11161, 
    11162, 
    11163, 
    11164, 
    11165, 
    11166, 
    11167, 
    11168, 
    11169, 
    11170, 
    11171, 
    11172, 
    11173, 
    11174, 
    11175, 
    11176, 
    11177, 
    11178, 
    11179, 
    11180, 
    11181, 
    11182, 
    11183, 
    11184, 
    11185, 
    11186, 
    11187, 
    11188, 
    11189, 
    11190, 
    11191, 
    11192, 
    11193, 
    11194, 
    11195, 
    11196, 
    11197, 
    11198, 
    11199, 
    11200, 
    11201, 
    11202, 
    11203, 
    11204, 
    11205, 
    11206, 
    11207, 
    11208, 
    11209, 
    11210, 
    11211, 
    11212, 
    11213, 
    11214, 
    11215, 
    11216, 
    11217, 
    11218, 
    11219, 
    11220, 
    11221, 
    11222, 
    11223, 
    11224, 
    11225, 
    11226, 
    11227, 
    11228, 
    11229, 
    11230, 
    11231, 
    11232, 
    11233, 
    11234, 
    11235, 
    11236, 
    11237, 
    11238, 
    11239, 
    11240, 
    11241, 
    11242, 
    11243, 
    11244, 
    11245, 
    11246, 
    11247, 
    11248, 
    11249, 
    11250, 
    11251, 
    11252, 
    11253, 
    11254, 
    11255, 
    11256, 
    11257, 
    11258, 
    11259, 
    11260, 
    11261, 
    11262, 
    11263, 
    11264, 
    11265, 
    11266, 
    11267, 
    11268, 
    11269, 
    11270, 
    11271, 
    11272, 
    11273, 
    11274, 
    11275, 
    11276, 
    11277, 
    11278, 
    11279, 
    11280, 
    11281, 
    11282, 
    11283, 
    11284, 
    11285, 
    11286, 
    11287, 
    11288, 
    11289, 
    11290, 
    11291, 
    11292, 
    11293, 
    11294, 
    11295, 
    11296, 
    11297, 
    11298, 
    11299, 
    11300, 
    11301, 
    11302, 
    11303, 
    11304, 
    11305, 
    11306, 
    11307, 
    11308, 
    11309, 
    11310, 
    11311, 
    11312, 
    11313, 
    11314, 
    11315, 
    11316, 
    11317, 
    11318, 
    11319, 
    11320, 
    11321, 
    11322, 
    11323, 
    11324, 
    11325, 
    11326, 
    11327, 
    11328, 
    11329, 
    11330, 
    11331, 
    11332, 
    11333, 
    11334, 
    11335, 
    11336, 
    11337, 
    11338, 
    11339, 
    11340, 
    11341, 
    11342, 
    11343, 
    11344, 
    11345, 
    11346, 
    11347, 
    11348, 
    11349, 
    11350, 
    11351, 
    11352, 
    11353, 
    11354, 
    11355, 
    11356, 
    11357, 
    11358, 
    11359, 
    11360, 
    11361, 
    11362, 
    11363, 
    11364, 
    11365, 
    11366, 
    11367, 
    11368, 
    11369, 
    11370, 
    11371, 
    11372, 
    11373, 
    11374, 
    11375, 
    11376, 
    11377, 
    11378, 
    11379, 
    11380, 
    11381, 
    11382, 
    11383, 
    11384, 
    11385, 
    11386, 
    11387, 
    11388, 
    11389, 
    11390, 
    11391, 
    11392, 
    11393, 
    11394, 
    11395, 
    11396, 
    11397, 
    11398, 
    11399, 
    11400, 
    11401, 
    11402, 
    11403, 
    11404, 
    11405, 
    11406, 
    11407, 
    11408, 
    11409, 
    11410, 
    11411, 
    11412, 
    11413, 
    11414, 
    11415, 
    11416, 
    11417, 
    11418, 
    11419, 
    11420, 
    11421, 
    11422, 
    11423, 
    11424, 
    11425, 
    11426, 
    11427, 
    11428, 
    11429, 
    11430, 
    11431, 
    11432, 
    11433, 
    11434, 
    11435, 
    11436, 
    11437, 
    11438, 
    11439, 
    11440, 
    11441, 
    11442, 
    11443, 
    11444, 
    11445, 
    11446, 
    11447, 
    11448, 
    11449, 
    11450, 
    11451, 
    11452, 
    11453, 
    11454, 
    11455, 
    11456, 
    11457, 
    11458, 
    11459, 
    11460, 
    11461, 
    11462, 
    11463, 
    11464, 
    11465, 
    11466, 
    11467, 
    11468, 
    11469, 
    11470, 
    11471, 
    11472, 
    11473, 
    11474, 
    11475, 
    11476, 
    11477, 
    11478, 
    11479, 
    11480, 
    11481, 
    11482, 
    11483, 
    11484, 
    11485, 
    11486, 
    11487, 
    11488, 
    11489, 
    11490, 
    11491, 
    11492, 
    11493, 
    11494, 
    11495, 
    11496, 
    11497, 
    11498, 
    11499, 
    11500, 
    11501, 
    11502, 
    11503, 
    11504, 
    11505, 
    11506, 
    11507, 
    11508, 
    11509, 
    11510, 
    11511, 
    11512, 
    11513, 
    11514, 
    11515, 
    11516, 
    11517, 
    11518, 
    11519, 
    11520, 
    11521, 
    11522, 
    11523, 
    11524, 
    11525, 
    11526, 
    11527, 
    11528, 
    11529, 
    11530, 
    11531, 
    11532, 
    11533, 
    11534, 
    11535, 
    11536, 
    11537, 
    11538, 
    11539, 
    11540, 
    11541, 
    11542, 
    11543, 
    11544, 
    11545, 
    11546, 
    11547, 
    11548, 
    11549, 
    11550, 
    11551, 
    11552, 
    11553, 
    11554, 
    11555, 
    11556, 
    11557, 
    11558, 
    11559, 
    11560, 
    11561, 
    11562, 
    11563, 
    11564, 
    11565, 
    11566, 
    11567, 
    11568, 
    11569, 
    11570, 
    11571, 
    11572, 
    11573, 
    11574, 
    11575, 
    11576, 
    11577, 
    11578, 
    11579, 
    11580, 
    11581, 
    11582, 
    11583, 
    11584, 
    11585, 
    11586, 
    11587, 
    11588, 
    11589, 
    11590, 
    11591, 
    11592, 
    11593, 
    11594, 
    11595, 
    11596, 
    11597, 
    11598, 
    11599, 
    11600, 
    11601, 
    11602, 
    11603, 
    11604, 
    11605, 
    11606, 
    11607, 
    11608, 
    11609, 
    11610, 
    11611, 
    11612, 
    11613, 
    11614, 
    11615, 
    11616, 
    11617, 
    11618, 
    11619, 
    11620, 
    11621, 
    11622, 
    11623, 
    11624, 
    11625, 
    11626, 
    11627, 
    11628, 
    11629, 
    11630, 
    11631, 
    11632, 
    11633, 
    11634, 
    11635, 
    11636, 
    11637, 
    11638, 
    11639, 
    11640, 
    11641, 
    11642, 
    11643, 
    11644, 
    11645, 
    11646, 
    11647, 
    11648, 
    11649, 
    11650, 
    11651, 
    11652, 
    11653, 
    11654, 
    11655, 
    11656, 
    11657, 
    11658, 
    11659, 
    11660, 
    11661, 
    11662, 
    11663, 
    11664, 
    11665, 
    11666, 
    11667, 
    11668, 
    11669, 
    11670, 
    11671, 
    11672, 
    11673, 
    11674, 
    11675, 
    11676, 
    11677, 
    11678, 
    11679, 
    11680, 
    11681, 
    11682, 
    11683, 
    11684, 
    11685, 
    11686, 
    11687, 
    11688, 
    11689, 
    11690, 
    11691, 
    11692, 
    11693, 
    11694, 
    11695, 
    11696, 
    11697, 
    11698, 
    11699, 
    11700, 
    11701, 
    11702, 
    11703, 
    11704, 
    11705, 
    11706, 
    11707, 
    11708, 
    11709, 
    11710, 
    11711, 
    11712, 
    11713, 
    11714, 
    11715, 
    11716, 
    11717, 
    11718, 
    11719, 
    11720, 
    11721, 
    11722, 
    11723, 
    11724, 
    11725, 
    11726, 
    11727, 
    11728, 
    11729, 
    11730, 
    11731, 
    11732, 
    11733, 
    11734, 
    11735, 
    11736, 
    11737, 
    11738, 
    11739, 
    11740, 
    11741, 
    11742, 
    11743, 
    11744, 
    11745, 
    11746, 
    11747, 
    11748, 
    11749, 
    11750, 
    11751, 
    11752, 
    11753, 
    11754, 
    11755, 
    11756, 
    11757, 
    11758, 
    11759, 
    11760, 
    11761, 
    11762, 
    11763, 
    11764, 
    11765, 
    11766, 
    11767, 
    11768, 
    11769, 
    11770, 
    11771, 
    11772, 
    11773, 
    11774, 
    11775, 
    11776, 
    11777, 
    11778, 
    11779, 
    11780, 
    11781, 
    11782, 
    11783, 
    11784, 
    11785, 
    11786, 
    11787, 
    11788, 
    11789, 
    11790, 
    11791, 
    11792, 
    11793, 
    11794, 
    11795, 
    11796, 
    11797, 
    11798, 
    11799, 
    11800, 
    11801, 
    11802, 
    11803, 
    11804, 
    11805, 
    11806, 
    11807, 
    11808, 
    11809, 
    11810, 
    11811, 
    11812, 
    11813, 
    11814, 
    11815, 
    11816, 
    11817, 
    11818, 
    11819, 
    11820, 
    11821, 
    11822, 
    11823, 
    11824, 
    11825, 
    11826, 
    11827, 
    11828, 
    11829, 
    11830, 
    11831, 
    11832, 
    11833, 
    11834, 
    11835, 
    11836, 
    11837, 
    11838, 
    11839, 
    11840, 
    11841, 
    11842, 
    11843, 
    11844, 
    11845, 
    11846, 
    11847, 
    11848, 
    11849, 
    11850, 
    11851, 
    11852, 
    11853, 
    11854, 
    11855, 
    11856, 
    11857, 
    11858, 
    11859, 
    11860, 
    11861, 
    11862, 
    11863, 
    11864, 
    11865, 
    11866, 
    11867, 
    11868, 
    11869, 
    11870, 
    11871, 
    11872, 
    11873, 
    11874, 
    11875, 
    11876, 
    11877, 
    11878, 
    11879, 
    11880, 
    11881, 
    11882, 
    11883, 
    11884, 
    11885, 
    11886, 
    11887, 
    11888, 
    11889, 
    11890, 
    11891, 
    11892, 
    11893, 
    11894, 
    11895, 
    11896, 
    11897, 
    11898, 
    11899, 
    11900, 
    11901, 
    11902, 
    11903, 
    11904, 
    11905, 
    11906, 
    11907, 
    11908, 
    11909, 
    11910, 
    11911, 
    11912, 
    11913, 
    11914, 
    11915, 
    11916, 
    11917, 
    11918, 
    11919, 
    11920, 
    11921, 
    11922, 
    11923, 
    11924, 
    11925, 
    11926, 
    11927, 
    11928, 
    11929, 
    11930, 
    11931, 
    11932, 
    11933, 
    11934, 
    11935, 
    11936, 
    11937, 
    11938, 
    11939, 
    11940, 
    11941, 
    11942, 
    11943, 
    11944, 
    11945, 
    11946, 
    11947, 
    11948, 
    11949, 
    11950, 
    11951, 
    11952, 
    11953, 
    11954, 
    11955, 
    11956, 
    11957, 
    11958, 
    11959, 
    11960, 
    11961, 
    11962, 
    11963, 
    11964, 
    11965, 
    11966, 
    11967, 
    11968, 
    11969, 
    11970, 
    11971, 
    11972, 
    11973, 
    11974, 
    11975, 
    11976, 
    11977, 
    11978, 
    11979, 
    11980, 
    11981, 
    11982, 
    11983, 
    11984, 
    11985, 
    11986, 
    11987, 
    11988, 
    11989, 
    11990, 
    11991, 
    11992, 
    11993, 
    11994, 
    11995, 
    11996, 
    11997, 
    11998, 
    11999, 
    12000, 
    12001, 
    12002, 
    12003, 
    12004, 
    12005, 
    12006, 
    12007, 
    12008, 
    12009, 
    12010, 
    12011, 
    12012, 
    12013, 
    12014, 
    12015, 
    12016, 
    12017, 
    12018, 
    12019, 
    12020, 
    12021, 
    12022, 
    12023, 
    12024, 
    12025, 
    12026, 
    12027, 
    12028, 
    12029, 
    12030, 
    12031, 
    12032, 
    12033, 
    12034, 
    12035, 
    12036, 
    12037, 
    12038, 
    12039, 
    12040, 
    12041, 
    12042, 
    12043, 
    12044, 
    12045, 
    12046, 
    12047, 
    12048, 
    12049, 
    12050, 
    12051, 
    12052, 
    12053, 
    12054, 
    12055, 
    12056, 
    12057, 
    12058, 
    12059, 
    12060, 
    12061, 
    12062, 
    12063, 
    12064, 
    12065, 
    12066, 
    12067, 
    12068, 
    12069, 
    12070, 
    12071, 
    12072, 
    12073, 
    12074, 
    12075, 
    12076, 
    12077, 
    12078, 
    12079, 
    12080, 
    12081, 
    12082, 
    12083, 
    12084, 
    12085, 
    12086, 
    12087, 
    12088, 
    12089, 
    12090, 
    12091, 
    12092, 
    12093, 
    12094, 
    12095, 
    12096, 
    12097, 
    12098, 
    12099, 
    12100, 
    12101, 
    12102, 
    12103, 
    12104, 
    12105, 
    12106, 
    12107, 
    12108, 
    12109, 
    12110, 
    12111, 
    12112, 
    12113, 
    12114, 
    12115, 
    12116, 
    12117, 
    12118, 
    12119, 
    12120, 
    12121, 
    12122, 
    12123, 
    12124, 
    12125, 
    12126, 
    12127, 
    12128, 
    12129, 
    12130, 
    12131, 
    12132, 
    12133, 
    12134, 
    12135, 
    12136, 
    12137, 
    12138, 
    12139, 
    12140, 
    12141, 
    12142, 
    12143, 
    12144, 
    12145, 
    12146, 
    12147, 
    12148, 
    12149, 
    12150, 
    12151, 
    12152, 
    12153, 
    12154, 
    12155, 
    12156, 
    12157, 
    12158, 
    12159, 
    12160, 
    12161, 
    12162, 
    12163, 
    12164, 
    12165, 
    12166, 
    12167, 
    12168, 
    12169, 
    12170, 
    12171, 
    12172, 
    12173, 
    12174, 
    12175, 
    12176, 
    12177, 
    12178, 
    12179, 
    12180, 
    12181, 
    12182, 
    12183, 
    12184, 
    12185, 
    12186, 
    12187, 
    12188, 
    12189, 
    12190, 
    12191, 
    12192, 
    12193, 
    12194, 
    12195, 
    12196, 
    12197, 
    12198, 
    12199, 
    12200, 
    12201, 
    12202, 
    12203, 
    12204, 
    12205, 
    12206, 
    12207, 
    12208, 
    12209, 
    12210, 
    12211, 
    12212, 
    12213, 
    12214, 
    12215, 
    12216, 
    12217, 
    12218, 
    12219, 
    12220, 
    12221, 
    12222, 
    12223, 
    12224, 
    12225, 
    12226, 
    12227, 
    12228, 
    12229, 
    12230, 
    12231, 
    12232, 
    12233, 
    12234, 
    12235, 
    12236, 
    12237, 
    12238, 
    12239, 
    12240, 
    12241, 
    12242, 
    12243, 
    12244, 
    12245, 
    12246, 
    12247, 
    12248, 
    12249, 
    12250, 
    12251, 
    12252, 
    12253, 
    12254, 
    12255, 
    12256, 
    12257, 
    12258, 
    12259, 
    12260, 
    12261, 
    12262, 
    12263, 
    12264, 
    12265, 
    12266, 
    12267, 
    12268, 
    12269, 
    12270, 
    12271, 
    12272, 
    12273, 
    12274, 
    12275, 
    12276, 
    12277, 
    12278, 
    12279, 
    12280, 
    12281, 
    12282, 
    12283, 
    12284, 
    12285, 
    12286, 
    12287, 
    12288, 
    12289, 
    12290, 
    12291, 
    12292, 
    12293, 
    12294, 
    12295, 
    12296, 
    12297, 
    12298, 
    12299, 
    12300, 
    12301, 
    12302, 
    12303, 
    12304, 
    12305, 
    12306, 
    12307, 
    12308, 
    12309, 
    12310, 
    12311, 
    12312, 
    12313, 
    12314, 
    12315, 
    12316, 
    12317, 
    12318, 
    12319, 
    12320, 
    12321, 
    12322, 
    12323, 
    12324, 
    12325, 
    12326, 
    12327, 
    12328, 
    12329, 
    12330, 
    12331, 
    12332, 
    12333, 
    12334, 
    12335, 
    12336, 
    12337, 
    12338, 
    12339, 
    12340, 
    12341, 
    12342, 
    12343, 
    12344, 
    12345, 
    12346, 
    12347, 
    12348, 
    12349, 
    12350, 
    12351, 
    12352, 
    12353, 
    12354, 
    12355, 
    12356, 
    12357, 
    12358, 
    12359, 
    12360, 
    12361, 
    12362, 
    12363, 
    12364, 
    12365, 
    12366, 
    12367, 
    12368, 
    12369, 
    12370, 
    12371, 
    12372, 
    12373, 
    12374, 
    12375, 
    12376, 
    12377, 
    12378, 
    12379, 
    12380, 
    12381, 
    12382, 
    12383, 
    12384, 
    12385, 
    12386, 
    12387, 
    12388, 
    12389, 
    12390, 
    12391, 
    12392, 
    12393, 
    12394, 
    12395, 
    12396, 
    12397, 
    12398, 
    12399, 
    12400, 
    12401, 
    12402, 
    12403, 
    12404, 
    12405, 
    12406, 
    12407, 
    12408, 
    12409, 
    12410, 
    12411, 
    12412, 
    12413, 
    12414, 
    12415, 
    12416, 
    12417, 
    12418, 
    12419, 
    12420, 
    12421, 
    12422, 
    12423, 
    12424, 
    12425, 
    12426, 
    12427, 
    12428, 
    12429, 
    12430, 
    12431, 
    12432, 
    12433, 
    12434, 
    12435, 
    12436, 
    12437, 
    12438, 
    12439, 
    12440, 
    12441, 
    12442, 
    12443, 
    12444, 
    12445, 
    12446, 
    12447, 
    12448, 
    12449, 
    12450, 
    12451, 
    12452, 
    12453, 
    12454, 
    12455, 
    12456, 
    12457, 
    12458, 
    12459, 
    12460, 
    12461, 
    12462, 
    12463, 
    12464, 
    12465, 
    12466, 
    12467, 
    12468, 
    12469, 
    12470, 
    12471, 
    12472, 
    12473, 
    12474, 
    12475, 
    12476, 
    12477, 
    12478, 
    12479, 
    12480, 
    12481, 
    12482, 
    12483, 
    12484, 
    12485, 
    12486, 
    12487, 
    12488, 
    12489, 
    12490, 
    12491, 
    12492, 
    12493, 
    12494, 
    12495, 
    12496, 
    12497, 
    12498, 
    12499, 
    12500, 
    12501, 
    12502, 
    12503, 
    12504, 
    12505, 
    12506, 
    12507, 
    12508, 
    12509, 
    12510, 
    12511, 
    12512, 
    12513, 
    12514, 
    12515, 
    12516, 
    12517, 
    12518, 
    12519, 
    12520, 
    12521, 
    12522, 
    12523, 
    12524, 
    12525, 
    12526, 
    12527, 
    12528, 
    12529, 
    12530, 
    12531, 
    12532, 
    12533, 
    12534, 
    12535, 
    12536, 
    12537, 
    12538, 
    12539, 
    12540, 
    12541, 
    12542, 
    12543, 
    12544, 
    12545, 
    12546, 
    12547, 
    12548, 
    12549, 
    12550, 
    12551, 
    12552, 
    12553, 
    12554, 
    12555, 
    12556, 
    12557, 
    12558, 
    12559, 
    12560, 
    12561, 
    12562, 
    12563, 
    12564, 
    12565, 
    12566, 
    12567, 
    12568, 
    12569, 
    12570, 
    12571, 
    12572, 
    12573, 
    12574, 
    12575, 
    12576, 
    12577, 
    12578, 
    12579, 
    12580, 
    12581, 
    12582, 
    12583, 
    12584, 
    12585, 
    12586, 
    12587, 
    12588, 
    12589, 
    12590, 
    12591, 
    12592, 
    12593, 
    12594, 
    12595, 
    12596, 
    12597, 
    12598, 
    12599, 
    12600, 
    12601, 
    12602, 
    12603, 
    12604, 
    12605, 
    12606, 
    12607, 
    12608, 
    12609, 
    12610, 
    12611, 
    12612, 
    12613, 
    12614, 
    12615, 
    12616, 
    12617, 
    12618, 
    12619, 
    12620, 
    12621, 
    12622, 
    12623, 
    12624, 
    12625, 
    12626, 
    12627, 
    12628, 
    12629, 
    12630, 
    12631, 
    12632, 
    12633, 
    12634, 
    12635, 
    12636, 
    12637, 
    12638, 
    12639, 
    12640, 
    12641, 
    12642, 
    12643, 
    12644, 
    12645, 
    12646, 
    12647, 
    12648, 
    12649, 
    12650, 
    12651, 
    12652, 
    12653, 
    12654, 
    12655, 
    12656, 
    12657, 
    12658, 
    12659, 
    12660, 
    12661, 
    12662, 
    12663, 
    12664, 
    12665, 
    12666, 
    12667, 
    12668, 
    12669, 
    12670, 
    12671, 
    12672, 
    12673, 
    12674, 
    12675, 
    12676, 
    12677, 
    12678, 
    12679, 
    12680, 
    12681, 
    12682, 
    12683, 
    12684, 
    12685, 
    12686, 
    12687, 
    12688, 
    12689, 
    12690, 
    12691, 
    12692, 
    12693, 
    12694, 
    12695, 
    12696, 
    12697, 
    12698, 
    12699, 
    12700, 
    12701, 
    12702, 
    12703, 
    12704, 
    12705, 
    12706, 
    12707, 
    12708, 
    12709, 
    12710, 
    12711, 
    12712, 
    12713, 
    12714, 
    12715, 
    12716, 
    12717, 
    12718, 
    12719, 
    12720, 
    12721, 
    12722, 
    12723, 
    12724, 
    12725, 
    12726, 
    12727, 
    12728, 
    12729, 
    12730, 
    12731, 
    12732, 
    12733, 
    12734, 
    12735, 
    12736, 
    12737, 
    12738, 
    12739, 
    12740, 
    12741, 
    12742, 
    12743, 
    12744, 
    12745, 
    12746, 
    12747, 
    12748, 
    12749, 
    12750, 
    12751 ;

 grid.cells.vertex_refs = 
    3693, 
    4860, 
    3398, 
    1741, 
    1628, 
    997, 
    190, 
    1741, 
    191, 
    6652, 
    187, 
    1968, 
    189, 
    6652, 
    1968, 
    189, 
    188, 
    6652, 
    3409, 
    982, 
    3080, 
    3961, 
    997, 
    1628, 
    3409, 
    4408, 
    3706, 
    6374, 
    3066, 
    3398, 
    4860, 
    6374, 
    3398, 
    5933, 
    6179, 
    6374, 
    799, 
    184, 
    2704, 
    1741, 
    189, 
    1968, 
    5775, 
    666, 
    183, 
    1457, 
    5775, 
    183, 
    4531, 
    1479, 
    5775, 
    5775, 
    1479, 
    666, 
    2090, 
    4864, 
    5027, 
    4705, 
    3238, 
    4531, 
    5066, 
    3071, 
    5582, 
    1626, 
    5066, 
    3549, 
    1626, 
    1037, 
    5503, 
    1041, 
    1479, 
    4531, 
    1041, 
    1214, 
    1479, 
    3080, 
    982, 
    1214, 
    5357, 
    3080, 
    838, 
    1310, 
    6392, 
    838, 
    2687, 
    5986, 
    5357, 
    3409, 
    3706, 
    5005, 
    5357, 
    5986, 
    3080, 
    6179, 
    5799, 
    4192, 
    4860, 
    5933, 
    6374, 
    4860, 
    6235, 
    5933, 
    5005, 
    609, 
    183, 
    1741, 
    190, 
    189, 
    187, 
    6652, 
    188, 
    1628, 
    1968, 
    185, 
    2704, 
    5645, 
    799, 
    997, 
    5762, 
    1741, 
    799, 
    1628, 
    185, 
    1968, 
    187, 
    186, 
    185, 
    1968, 
    186, 
    1628, 
    1741, 
    1968, 
    185, 
    184, 
    799, 
    666, 
    5005, 
    183, 
    2870, 
    5305, 
    1060, 
    1011, 
    3116, 
    2452, 
    3996, 
    1552, 
    2144, 
    5125, 
    4843, 
    3996, 
    3116, 
    5125, 
    2750, 
    4493, 
    2444, 
    5125, 
    4843, 
    3098, 
    4066, 
    3720, 
    1060, 
    3429, 
    670, 
    3720, 
    3429, 
    1529, 
    1132, 
    3720, 
    3720, 
    1132, 
    1817, 
    2483, 
    2899, 
    3427, 
    1132, 
    6310, 
    1027, 
    4141, 
    817, 
    2012, 
    4801, 
    4141, 
    2012, 
    1338, 
    4801, 
    2012, 
    2913, 
    5529, 
    4801, 
    5507, 
    3849, 
    1643, 
    3886, 
    5507, 
    4141, 
    3886, 
    2039, 
    5507, 
    4801, 
    3886, 
    4141, 
    1385, 
    2039, 
    3886, 
    3255, 
    2913, 
    4801, 
    2322, 
    3255, 
    1338, 
    2322, 
    1785, 
    3985, 
    2913, 
    1817, 
    2349, 
    1385, 
    5529, 
    2349, 
    3255, 
    3985, 
    4982, 
    1060, 
    3720, 
    1817, 
    1615, 
    781, 
    2039, 
    4350, 
    1615, 
    1385, 
    1027, 
    2767, 
    5450, 
    2349, 
    4350, 
    1385, 
    3482, 
    761, 
    3821, 
    4796, 
    1982, 
    3482, 
    4135, 
    1443, 
    2383, 
    3874, 
    4135, 
    2473, 
    3874, 
    1291, 
    6212, 
    4796, 
    1291, 
    1982, 
    2420, 
    4796, 
    1507, 
    2420, 
    1914, 
    4796, 
    1785, 
    1914, 
    1011, 
    3565, 
    1746, 
    2456, 
    1914, 
    3565, 
    2456, 
    1196, 
    2224, 
    4543, 
    1443, 
    5307, 
    2079, 
    4754, 
    939, 
    2079, 
    1746, 
    4754, 
    1192, 
    3872, 
    939, 
    4754, 
    5307, 
    4754, 
    2079, 
    3874, 
    6212, 
    4135, 
    1192, 
    4754, 
    5307, 
    5859, 
    1366, 
    1969, 
    1465, 
    5859, 
    2735, 
    1465, 
    1366, 
    5859, 
    5182, 
    1166, 
    1896, 
    5282, 
    5182, 
    2606, 
    1122, 
    5282, 
    2606, 
    1866, 
    2383, 
    5549, 
    6191, 
    3009, 
    2622, 
    5282, 
    6079, 
    5182, 
    5549, 
    3344, 
    6079, 
    1157, 
    310, 
    625, 
    4666, 
    1157, 
    625, 
    309, 
    4666, 
    625, 
    1045, 
    1806, 
    5104, 
    928, 
    2199, 
    1157, 
    2949, 
    3086, 
    3413, 
    4646, 
    1122, 
    2180, 
    1781, 
    4465, 
    3086, 
    4465, 
    6209, 
    5240, 
    5392, 
    1896, 
    2408, 
    4615, 
    5392, 
    2408, 
    2606, 
    5182, 
    5392, 
    1122, 
    2606, 
    2180, 
    1122, 
    1866, 
    5282, 
    2269, 
    983, 
    2103, 
    2022, 
    1722, 
    1358, 
    936, 
    1765, 
    1722, 
    1136, 
    172, 
    171, 
    6596, 
    174, 
    173, 
    1136, 
    173, 
    172, 
    788, 
    1735, 
    171, 
    901, 
    1701, 
    1136, 
    168, 
    788, 
    169, 
    170, 
    169, 
    788, 
    6092, 
    4496, 
    4846, 
    788, 
    6092, 
    4846, 
    3355, 
    4672, 
    6092, 
    1136, 
    1735, 
    901, 
    3355, 
    6092, 
    3022, 
    170, 
    788, 
    171, 
    3022, 
    167, 
    917, 
    171, 
    1735, 
    1136, 
    5759, 
    2797, 
    4757, 
    3191, 
    3361, 
    5838, 
    4771, 
    3760, 
    4025, 
    3689, 
    6507, 
    3392, 
    3472, 
    3760, 
    4603, 
    168, 
    167, 
    3022, 
    1703, 
    166, 
    165, 
    3014, 
    4839, 
    907, 
    1898, 
    166, 
    1703, 
    4839, 
    4664, 
    1703, 
    1169, 
    917, 
    1898, 
    4940, 
    917, 
    1169, 
    4672, 
    4496, 
    6092, 
    3191, 
    4672, 
    863, 
    3191, 
    2841, 
    4672, 
    3355, 
    917, 
    1811, 
    3355, 
    3022, 
    917, 
    863, 
    4672, 
    1811, 
    4846, 
    4289, 
    1735, 
    1811, 
    4672, 
    3355, 
    2841, 
    5465, 
    4496, 
    788, 
    168, 
    3022, 
    167, 
    166, 
    1898, 
    178, 
    4570, 
    1225, 
    175, 
    1701, 
    176, 
    3361, 
    1673, 
    715, 
    3361, 
    3191, 
    1673, 
    5955, 
    4025, 
    3662, 
    1922, 
    4251, 
    695, 
    1922, 
    4483, 
    4251, 
    3662, 
    5838, 
    3361, 
    715, 
    695, 
    5955, 
    6447, 
    5641, 
    5838, 
    5931, 
    6447, 
    5797, 
    5977, 
    5641, 
    6447, 
    5296, 
    5977, 
    5837, 
    5393, 
    5465, 
    5977, 
    4025, 
    3933, 
    3662, 
    3472, 
    3153, 
    6470, 
    2841, 
    4496, 
    4672, 
    5977, 
    6447, 
    5837, 
    2841, 
    5641, 
    5465, 
    3933, 
    4174, 
    5797, 
    4745, 
    5296, 
    2731, 
    1701, 
    901, 
    5393, 
    4846, 
    1735, 
    788, 
    3022, 
    6092, 
    788, 
    4496, 
    4289, 
    4846, 
    5465, 
    5641, 
    5977, 
    901, 
    1735, 
    4289, 
    3431, 
    682, 
    1323, 
    3102, 
    3431, 
    1323, 
    5759, 
    6470, 
    3153, 
    682, 
    4930, 
    4757, 
    3102, 
    2731, 
    5069, 
    1225, 
    3102, 
    1323, 
    3933, 
    6447, 
    5838, 
    6470, 
    6535, 
    5797, 
    3472, 
    6470, 
    4174, 
    6535, 
    5931, 
    5797, 
    5759, 
    6535, 
    6470, 
    5759, 
    4930, 
    6535, 
    5977, 
    5296, 
    5393, 
    5931, 
    5837, 
    6447, 
    5069, 
    2731, 
    5837, 
    1225, 
    4570, 
    3102, 
    5393, 
    901, 
    4289, 
    5465, 
    5393, 
    4289, 
    4496, 
    5465, 
    4289, 
    5838, 
    3662, 
    3933, 
    2841, 
    5838, 
    5641, 
    2841, 
    3191, 
    5838, 
    5296, 
    1701, 
    5393, 
    4940, 
    1169, 
    2210, 
    1978, 
    1017, 
    2119, 
    6698, 
    320, 
    319, 
    2086, 
    6698, 
    319, 
    629, 
    320, 
    6698, 
    629, 
    6698, 
    2086, 
    1539, 
    2086, 
    318, 
    2086, 
    630, 
    629, 
    318, 
    2086, 
    319, 
    1539, 
    686, 
    2086, 
    321, 
    1228, 
    322, 
    686, 
    321, 
    630, 
    4764, 
    317, 
    628, 
    4762, 
    4764, 
    628, 
    2133, 
    318, 
    4764, 
    5561, 
    1183, 
    3068, 
    4764, 
    4762, 
    2133, 
    316, 
    1183, 
    4762, 
    4762, 
    628, 
    316, 
    2216, 
    3068, 
    1183, 
    2381, 
    2216, 
    1183, 
    3491, 
    840, 
    2022, 
    4311, 
    5311, 
    3243, 
    4410, 
    840, 
    3491, 
    1539, 
    318, 
    2133, 
    4266, 
    2468, 
    4311, 
    2829, 
    4266, 
    2487, 
    2884, 
    2468, 
    4266, 
    1766, 
    2884, 
    4472, 
    1766, 
    985, 
    5488, 
    1440, 
    1655, 
    2216, 
    1440, 
    2077, 
    1655, 
    2381, 
    1440, 
    2216, 
    627, 
    2381, 
    1183, 
    784, 
    1440, 
    2381, 
    784, 
    973, 
    1440, 
    2086, 
    686, 
    630, 
    317, 
    4764, 
    318, 
    3068, 
    2216, 
    1655, 
    4410, 
    3068, 
    1655, 
    3243, 
    5311, 
    3491, 
    3401, 
    3068, 
    4410, 
    5311, 
    3401, 
    4410, 
    3491, 
    5311, 
    4410, 
    4311, 
    3696, 
    5311, 
    3963, 
    3696, 
    2468, 
    2884, 
    5488, 
    2468, 
    4513, 
    3871, 
    3602, 
    5922, 
    4513, 
    4313, 
    2691, 
    3871, 
    4513, 
    4313, 
    3602, 
    3295, 
    6489, 
    5922, 
    4313, 
    5260, 
    6489, 
    4096, 
    5260, 
    5737, 
    6489, 
    3963, 
    2691, 
    4513, 
    4096, 
    4313, 
    3295, 
    5561, 
    4762, 
    1183, 
    3401, 
    5561, 
    3068, 
    5737, 
    5260, 
    5561, 
    3401, 
    5737, 
    5561, 
    3401, 
    3696, 
    5737, 
    1228, 
    321, 
    686, 
    3295, 
    1228, 
    686, 
    323, 
    322, 
    1228, 
    2205, 
    154, 
    605, 
    3810, 
    1694, 
    1010, 
    153, 
    3768, 
    1642, 
    894, 
    1694, 
    3768, 
    604, 
    1337, 
    5455, 
    5455, 
    894, 
    3768, 
    151, 
    1337, 
    604, 
    5802, 
    6473, 
    4972, 
    5129, 
    4582, 
    6243, 
    5455, 
    1337, 
    894, 
    153, 
    5455, 
    3768, 
    152, 
    604, 
    5455, 
    2357, 
    603, 
    149, 
    6504, 
    1271, 
    1861, 
    4647, 
    6504, 
    1861, 
    6221, 
    5959, 
    6504, 
    4819, 
    5959, 
    5334, 
    1435, 
    1271, 
    6504, 
    151, 
    150, 
    1401, 
    1211, 
    159, 
    158, 
    157, 
    156, 
    1927, 
    1927, 
    905, 
    2031, 
    157, 
    1927, 
    158, 
    156, 
    905, 
    1927, 
    1642, 
    2205, 
    605, 
    1211, 
    1927, 
    2031, 
    156, 
    155, 
    905, 
    1667, 
    160, 
    857, 
    1211, 
    160, 
    159, 
    1927, 
    1211, 
    158, 
    857, 
    160, 
    1211, 
    2115, 
    1231, 
    1510, 
    1916, 
    4967, 
    3983, 
    857, 
    2422, 
    1667, 
    4967, 
    1542, 
    3983, 
    2422, 
    4967, 
    1916, 
    690, 
    1542, 
    4967, 
    1667, 
    161, 
    160, 
    2422, 
    1916, 
    1667, 
    2031, 
    2422, 
    857, 
    1510, 
    1941, 
    2422, 
    1199, 
    606, 
    1667, 
    4499, 
    3810, 
    1010, 
    155, 
    4499, 
    3656, 
    2205, 
    3810, 
    4499, 
    154, 
    2205, 
    155, 
    4499, 
    1010, 
    2115, 
    1642, 
    3810, 
    2205, 
    1642, 
    3768, 
    3810, 
    153, 
    1642, 
    605, 
    153, 
    152, 
    5455, 
    163, 
    6597, 
    164, 
    4425, 
    607, 
    162, 
    1703, 
    967, 
    907, 
    5134, 
    607, 
    1044, 
    1751, 
    967, 
    1044, 
    1199, 
    162, 
    606, 
    161, 
    1667, 
    606, 
    3983, 
    2135, 
    4425, 
    1916, 
    3983, 
    1199, 
    1542, 
    2135, 
    3983, 
    1667, 
    1916, 
    1199, 
    4813, 
    1296, 
    4004, 
    690, 
    4813, 
    1542, 
    690, 
    2721, 
    6188, 
    603, 
    1401, 
    150, 
    149, 
    887, 
    1834, 
    147, 
    887, 
    148, 
    144, 
    143, 
    6573, 
    6573, 
    909, 
    145, 
    144, 
    6573, 
    145, 
    143, 
    909, 
    6573, 
    909, 
    147, 
    146, 
    145, 
    909, 
    146, 
    143, 
    1224, 
    3797, 
    909, 
    887, 
    147, 
    729, 
    1568, 
    141, 
    1938, 
    1224, 
    143, 
    141, 
    1938, 
    142, 
    1568, 
    2156, 
    1938, 
    1261, 
    1568, 
    729, 
    1261, 
    1447, 
    2560, 
    148, 
    887, 
    149, 
    1568, 
    1938, 
    141, 
    2242, 
    1224, 
    2156, 
    1834, 
    2242, 
    1079, 
    887, 
    909, 
    2242, 
    143, 
    142, 
    1938, 
    140, 
    139, 
    729, 
    141, 
    140, 
    729, 
    685, 
    1279, 
    137, 
    4917, 
    2170, 
    1099, 
    6118, 
    4917, 
    3796, 
    4830, 
    2170, 
    4917, 
    3516, 
    6118, 
    3796, 
    4562, 
    1585, 
    4830, 
    4121, 
    1585, 
    751, 
    4917, 
    1099, 
    4054, 
    1256, 
    2170, 
    1585, 
    1256, 
    1099, 
    2170, 
    1131, 
    1256, 
    683, 
    1131, 
    1040, 
    2186, 
    2132, 
    1131, 
    683, 
    1040, 
    1803, 
    2186, 
    4912, 
    2641, 
    3787, 
    3764, 
    4912, 
    3787, 
    4029, 
    5055, 
    4912, 
    2744, 
    5093, 
    5447, 
    5055, 
    4273, 
    2641, 
    4255, 
    5055, 
    4029, 
    4255, 
    5187, 
    5055, 
    5447, 
    5365, 
    4029, 
    3764, 
    5447, 
    4029, 
    5093, 
    5224, 
    5447, 
    5187, 
    1120, 
    4481, 
    1861, 
    1271, 
    6003, 
    5179, 
    4983, 
    5928, 
    1577, 
    5129, 
    743, 
    1577, 
    1601, 
    5129, 
    1834, 
    5324, 
    2357, 
    1435, 
    5959, 
    2536, 
    6221, 
    4826, 
    5649, 
    5959, 
    6221, 
    5334, 
    4647, 
    4826, 
    6221, 
    3142, 
    1728, 
    932, 
    6050, 
    3142, 
    2783, 
    2626, 
    6050, 
    2783, 
    3013, 
    5627, 
    6050, 
    3013, 
    3348, 
    5627, 
    1634, 
    821, 
    807, 
    1891, 
    1165, 
    972, 
    4485, 
    1891, 
    972, 
    4485, 
    4276, 
    3155, 
    5111, 
    4485, 
    972, 
    5111, 
    5329, 
    4485, 
    1261, 
    729, 
    5091, 
    2786, 
    6146, 
    1279, 
    5916, 
    2670, 
    2786, 
    3018, 
    5916, 
    2631, 
    1891, 
    2670, 
    5916, 
    1472, 
    139, 
    6146, 
    3155, 
    1472, 
    1891, 
    6146, 
    1431, 
    1279, 
    1472, 
    6146, 
    2670, 
    139, 
    1431, 
    6146, 
    4471, 
    2794, 
    3151, 
    4741, 
    770, 
    1987, 
    807, 
    4741, 
    1987, 
    783, 
    2317, 
    5268, 
    3018, 
    1165, 
    5916, 
    5052, 
    3018, 
    2631, 
    2794, 
    5052, 
    2631, 
    2599, 
    2817, 
    5052, 
    1764, 
    1165, 
    3018, 
    2028, 
    4621, 
    4574, 
    1278, 
    1977, 
    4621, 
    1278, 
    862, 
    1977, 
    4506, 
    1059, 
    2143, 
    1981, 
    4506, 
    760, 
    1981, 
    5221, 
    4506, 
    5471, 
    4321, 
    4106, 
    4694, 
    5471, 
    4106, 
    4517, 
    4201, 
    5471, 
    1810, 
    4104, 
    3236, 
    2344, 
    1374, 
    4107, 
    2036, 
    3567, 
    1374, 
    3512, 
    3196, 
    3841, 
    3259, 
    1816, 
    5359, 
    2169, 
    1584, 
    2344, 
    1098, 
    2169, 
    1810, 
    1098, 
    4650, 
    5500, 
    5349, 
    3792, 
    862, 
    5636, 
    3554, 
    3241, 
    5349, 
    6446, 
    5630, 
    5793, 
    948, 
    1921, 
    6446, 
    5793, 
    5636, 
    5630, 
    6446, 
    5636, 
    1672, 
    2281, 
    6446, 
    1736, 
    948, 
    5793, 
    2644, 
    3031, 
    3196, 
    750, 
    2036, 
    1374, 
    2873, 
    2455, 
    6177, 
    3223, 
    2873, 
    2655, 
    5144, 
    5254, 
    2873, 
    6455, 
    2709, 
    2485, 
    4591, 
    6455, 
    5664, 
    6059, 
    2709, 
    6455, 
    4591, 
    5254, 
    6455, 
    5254, 
    5144, 
    6495, 
    2455, 
    5254, 
    4591, 
    5144, 
    6101, 
    6495, 
    3223, 
    5000, 
    5144, 
    5466, 
    2843, 
    3935, 
    3085, 
    5466, 
    5394, 
    5660, 
    2843, 
    5466, 
    3412, 
    5660, 
    5466, 
    3412, 
    3710, 
    5660, 
    3972, 
    4052, 
    3259, 
    4988, 
    2705, 
    2847, 
    3363, 
    5396, 
    4988, 
    5298, 
    4387, 
    3707, 
    5396, 
    5298, 
    3410, 
    3935, 
    4387, 
    5298, 
    5466, 
    3935, 
    3664, 
    2843, 
    3193, 
    4175, 
    5017, 
    3076, 
    3405, 
    5413, 
    5017, 
    4867, 
    3081, 
    5413, 
    4867, 
    3410, 
    2505, 
    5413, 
    5413, 
    5154, 
    5017, 
    4867, 
    5017, 
    3405, 
    5254, 
    6059, 
    6455, 
    4988, 
    3081, 
    2705, 
    3363, 
    4988, 
    2847, 
    3363, 
    3664, 
    5396, 
    5512, 
    6076, 
    3031, 
    5396, 
    3410, 
    3081, 
    4988, 
    5396, 
    3081, 
    3664, 
    5298, 
    5396, 
    6351, 
    3664, 
    3363, 
    6076, 
    6351, 
    3363, 
    5394, 
    5466, 
    6351, 
    4175, 
    3193, 
    3508, 
    4586, 
    4175, 
    3508, 
    3707, 
    4387, 
    3972, 
    3707, 
    3410, 
    5298, 
    3935, 
    2843, 
    4175, 
    3792, 
    2036, 
    862, 
    3512, 
    3792, 
    2648, 
    5843, 
    2648, 
    5630, 
    1588, 
    1790, 
    754, 
    6337, 
    3638, 
    5555, 
    6520, 
    6337, 
    4583, 
    5551, 
    3332, 
    6337, 
    1408, 
    2840, 
    3004, 
    1408, 
    1296, 
    2840, 
    4016, 
    3908, 
    3638, 
    4555, 
    1662, 
    2222, 
    1736, 
    4555, 
    2222, 
    2281, 
    3384, 
    4555, 
    6446, 
    2281, 
    1736, 
    1278, 
    3384, 
    2281, 
    4597, 
    1190, 
    2222, 
    6136, 
    4073, 
    4597, 
    2078, 
    6136, 
    937, 
    2078, 
    6018, 
    6136, 
    6018, 
    1441, 
    4714, 
    6136, 
    6018, 
    4073, 
    2078, 
    1441, 
    6018, 
    5011, 
    4611, 
    4857, 
    4744, 
    5011, 
    4857, 
    4916, 
    1723, 
    5011, 
    6018, 
    4714, 
    4073, 
    2995, 
    1865, 
    1120, 
    2179, 
    5336, 
    1120, 
    6007, 
    1501, 
    3754, 
    1921, 
    4030, 
    1452, 
    2111, 
    2995, 
    1003, 
    6007, 
    1865, 
    2995, 
    2111, 
    6007, 
    2995, 
    3754, 
    1865, 
    6007, 
    2417, 
    3754, 
    1501, 
    2382, 
    1865, 
    3754, 
    2417, 
    4714, 
    3754, 
    4815, 
    2417, 
    1501, 
    4714, 
    1441, 
    2382, 
    1910, 
    4714, 
    2417, 
    1910, 
    4073, 
    4714, 
    3253, 
    2078, 
    937, 
    4916, 
    3253, 
    937, 
    1723, 
    4916, 
    937, 
    4744, 
    3562, 
    4916, 
    4620, 
    4422, 
    3562, 
    3074, 
    4791, 
    2698, 
    3222, 
    4422, 
    4620, 
    3222, 
    3533, 
    4422, 
    4422, 
    3533, 
    4210, 
    3253, 
    4422, 
    4210, 
    3562, 
    2698, 
    4620, 
    2912, 
    2498, 
    2619, 
    2654, 
    2912, 
    1017, 
    2654, 
    4228, 
    2912, 
    4651, 
    4468, 
    4601, 
    2328, 
    4651, 
    4601, 
    1343, 
    2016, 
    5690, 
    5690, 
    4651, 
    1343, 
    4915, 
    5690, 
    2016, 
    4915, 
    5655, 
    6124, 
    825, 
    4915, 
    2016, 
    4743, 
    5655, 
    4915, 
    4939, 
    4770, 
    4260, 
    2836, 
    4939, 
    4260, 
    4002, 
    4228, 
    4939, 
    4743, 
    4915, 
    4482, 
    6352, 
    6162, 
    6263, 
    6357, 
    6358, 
    5811, 
    5691, 
    6340, 
    5623, 
    5501, 
    5975, 
    6380, 
    5655, 
    4743, 
    6204, 
    6124, 
    5690, 
    4915, 
    5976, 
    6124, 
    5655, 
    4468, 
    4651, 
    6124, 
    4482, 
    4274, 
    4743, 
    4743, 
    4274, 
    4568, 
    1649, 
    4482, 
    825, 
    1649, 
    4737, 
    4482, 
    4049, 
    4568, 
    4274, 
    2872, 
    3222, 
    4620, 
    2812, 
    2872, 
    2454, 
    3253, 
    4210, 
    2078, 
    5460, 
    5384, 
    3222, 
    2812, 
    5460, 
    2872, 
    5648, 
    5520, 
    3359, 
    5769, 
    5648, 
    5606, 
    5726, 
    5769, 
    5606, 
    5460, 
    2812, 
    5801, 
    6308, 
    5706, 
    5501, 
    5769, 
    5801, 
    5648, 
    2812, 
    5706, 
    5801, 
    3533, 
    3811, 
    4210, 
    5384, 
    5290, 
    3533, 
    2872, 
    5460, 
    3222, 
    5460, 
    5769, 
    5384, 
    4210, 
    1441, 
    2078, 
    3562, 
    4422, 
    3253, 
    3811, 
    1441, 
    4210, 
    5190, 
    6067, 
    4481, 
    2382, 
    1441, 
    3811, 
    5268, 
    4741, 
    783, 
    2071, 
    2741, 
    926, 
    3673, 
    2474, 
    3507, 
    6101, 
    3412, 
    3085, 
    6495, 
    6101, 
    3085, 
    6059, 
    6495, 
    3085, 
    6059, 
    5254, 
    6495, 
    5144, 
    5000, 
    6101, 
    6101, 
    4279, 
    3412, 
    3534, 
    5000, 
    3223, 
    3534, 
    5201, 
    5000, 
    4057, 
    3710, 
    4279, 
    4784, 
    3508, 
    4945, 
    4945, 
    2843, 
    3710, 
    3534, 
    2890, 
    3372, 
    3534, 
    3223, 
    2655, 
    5302, 
    3798, 
    6254, 
    3372, 
    5302, 
    5201, 
    3673, 
    3942, 
    5400, 
    4279, 
    3710, 
    3412, 
    5201, 
    4057, 
    5000, 
    3372, 
    5201, 
    3534, 
    6254, 
    4057, 
    5201, 
    5302, 
    6254, 
    5201, 
    3798, 
    4057, 
    6254, 
    3798, 
    3975, 
    4057, 
    3372, 
    3673, 
    5302, 
    4945, 
    3508, 
    3193, 
    4204, 
    4784, 
    3975, 
    4204, 
    4614, 
    4784, 
    3798, 
    4204, 
    3975, 
    3517, 
    3205, 
    4415, 
    3664, 
    6351, 
    5466, 
    5144, 
    2873, 
    3223, 
    4279, 
    6101, 
    5000, 
    3085, 
    2709, 
    6059, 
    2655, 
    2890, 
    3534, 
    3827, 
    3470, 
    1243, 
    3972, 
    2917, 
    3707, 
    6132, 
    1706, 
    912, 
    2741, 
    6132, 
    4602, 
    2741, 
    1706, 
    6132, 
    1243, 
    3205, 
    2257, 
    708, 
    4614, 
    1950, 
    3517, 
    3798, 
    5302, 
    4415, 
    4204, 
    3517, 
    1243, 
    4415, 
    3205, 
    1243, 
    1950, 
    4415, 
    4057, 
    4279, 
    5000, 
    2434, 
    2257, 
    3205, 
    2257, 
    2434, 
    1706, 
    2624, 
    1014, 
    1788, 
    4586, 
    3972, 
    4387, 
    2143, 
    4052, 
    4758, 
    2143, 
    1059, 
    4052, 
    5660, 
    3710, 
    2843, 
    4758, 
    4586, 
    3508, 
    2143, 
    4758, 
    1551, 
    4052, 
    4586, 
    4758, 
    4204, 
    3798, 
    3517, 
    4945, 
    3975, 
    4784, 
    2843, 
    4945, 
    3193, 
    3710, 
    3975, 
    4945, 
    3710, 
    4057, 
    3975, 
    3789, 
    708, 
    1551, 
    4784, 
    4614, 
    3789, 
    4614, 
    708, 
    3789, 
    3011, 
    4676, 
    2624, 
    5083, 
    1014, 
    1003, 
    1779, 
    5083, 
    1003, 
    1779, 
    1788, 
    5083, 
    1779, 
    1616, 
    1788, 
    5336, 
    2179, 
    4785, 
    2995, 
    5336, 
    1003, 
    2995, 
    1120, 
    5336, 
    2317, 
    1616, 
    1779, 
    4785, 
    2317, 
    1779, 
    5268, 
    770, 
    4741, 
    4785, 
    5268, 
    2317, 
    1605, 
    770, 
    5268, 
    6261, 
    2633, 
    3019, 
    1616, 
    6261, 
    3019, 
    783, 
    5553, 
    6261, 
    4512, 
    1099, 
    1961, 
    725, 
    4512, 
    1961, 
    1848, 
    1099, 
    4512, 
    3942, 
    3507, 
    3192, 
    2434, 
    5400, 
    3942, 
    3372, 
    2474, 
    3673, 
    5484, 
    821, 
    1634, 
    5484, 
    3170, 
    821, 
    1764, 
    5484, 
    1634, 
    1764, 
    3018, 
    6035, 
    6432, 
    5572, 
    5249, 
    5677, 
    6432, 
    5299, 
    5777, 
    5572, 
    6432, 
    2817, 
    5777, 
    5677, 
    2817, 
    2599, 
    5777, 
    6035, 
    2817, 
    5484, 
    1764, 
    6035, 
    5484, 
    3018, 
    5052, 
    6035, 
    5572, 
    2433, 
    5249, 
    5138, 
    4278, 
    2369, 
    1417, 
    5138, 
    2369, 
    4996, 
    5489, 
    5138, 
    3680, 
    4996, 
    2443, 
    4842, 
    5658, 
    4996, 
    3049, 
    4492, 
    4671, 
    4663, 
    3796, 
    4487, 
    5553, 
    783, 
    1993, 
    821, 
    6245, 
    1993, 
    5200, 
    2633, 
    5553, 
    5586, 
    3011, 
    2624, 
    5200, 
    5720, 
    5728, 
    3345, 
    3011, 
    5586, 
    6458, 
    5519, 
    5679, 
    6458, 
    5720, 
    5519, 
    5849, 
    6458, 
    5679, 
    5861, 
    5720, 
    6458, 
    5985, 
    5998, 
    5849, 
    5728, 
    5720, 
    5861, 
    2633, 
    5728, 
    5586, 
    2633, 
    5200, 
    5728, 
    5200, 
    5299, 
    5720, 
    4166, 
    3822, 
    4088, 
    5510, 
    2455, 
    4591, 
    5510, 
    3822, 
    6177, 
    6307, 
    4088, 
    5510, 
    5925, 
    4507, 
    4303, 
    3041, 
    5925, 
    2657, 
    6525, 
    5633, 
    4687, 
    3041, 
    6525, 
    5925, 
    3041, 
    5633, 
    6525, 
    3649, 
    3919, 
    4303, 
    3919, 
    4166, 
    4088, 
    5861, 
    5586, 
    5728, 
    3516, 
    6386, 
    3202, 
    6177, 
    2455, 
    5510, 
    3546, 
    6177, 
    3822, 
    3546, 
    2655, 
    6177, 
    5946, 
    6379, 
    6386, 
    2655, 
    2873, 
    6177, 
    4303, 
    3919, 
    4088, 
    6261, 
    1616, 
    783, 
    5586, 
    3019, 
    2633, 
    2624, 
    1788, 
    3019, 
    5083, 
    1788, 
    1014, 
    5963, 
    5299, 
    5200, 
    6245, 
    5677, 
    5963, 
    1993, 
    6245, 
    5553, 
    821, 
    3170, 
    6245, 
    3170, 
    2817, 
    5677, 
    4125, 
    5303, 
    3217, 
    5266, 
    4125, 
    3861, 
    5166, 
    5266, 
    3861, 
    3553, 
    3240, 
    5266, 
    5303, 
    2448, 
    2866, 
    5364, 
    4334, 
    4125, 
    2738, 
    1572, 
    5404, 
    2484, 
    1967, 
    736, 
    4125, 
    3217, 
    3861, 
    4791, 
    2454, 
    2872, 
    4791, 
    2758, 
    2454, 
    2698, 
    4791, 
    4620, 
    3074, 
    2758, 
    4791, 
    5011, 
    2270, 
    4611, 
    5016, 
    3006, 
    2498, 
    4863, 
    3647, 
    3342, 
    3123, 
    4692, 
    3449, 
    3701, 
    3647, 
    4692, 
    3123, 
    5508, 
    4692, 
    5603, 
    4155, 
    6295, 
    3553, 
    6189, 
    3240, 
    4569, 
    3074, 
    2698, 
    4563, 
    4508, 
    5698, 
    4305, 
    5708, 
    4508, 
    6025, 
    4305, 
    4091, 
    3403, 
    3074, 
    5128, 
    2758, 
    3403, 
    5508, 
    4744, 
    2698, 
    3562, 
    4366, 
    4689, 
    4782, 
    4689, 
    5128, 
    4569, 
    2479, 
    3006, 
    3342, 
    4228, 
    2498, 
    2912, 
    4601, 
    4770, 
    2654, 
    4002, 
    2498, 
    4228, 
    5502, 
    4002, 
    4939, 
    3186, 
    5502, 
    2836, 
    3737, 
    4002, 
    5502, 
    3737, 
    4863, 
    5016, 
    5884, 
    3449, 
    3737, 
    3186, 
    5884, 
    5502, 
    3186, 
    5306, 
    5884, 
    3449, 
    4692, 
    4863, 
    4738, 
    4091, 
    4305, 
    6189, 
    6082, 
    4738, 
    4366, 
    6522, 
    4563, 
    3553, 
    6082, 
    6189, 
    6367, 
    4092, 
    5842, 
    6484, 
    6367, 
    5842, 
    6082, 
    3826, 
    6367, 
    2479, 
    2895, 
    3006, 
    5896, 
    2270, 
    3682, 
    5458, 
    5896, 
    3682, 
    2993, 
    1266, 
    5896, 
    2460, 
    2993, 
    2603, 
    1266, 
    2270, 
    5896, 
    2484, 
    3906, 
    1967, 
    1967, 
    3906, 
    1266, 
    4397, 
    937, 
    6136, 
    3682, 
    4397, 
    3385, 
    1723, 
    937, 
    4397, 
    4073, 
    1190, 
    4597, 
    5458, 
    848, 
    2028, 
    2993, 
    5458, 
    2603, 
    3385, 
    848, 
    5458, 
    3682, 
    3385, 
    5458, 
    1723, 
    3682, 
    2270, 
    1723, 
    4397, 
    3682, 
    1662, 
    848, 
    3385, 
    2603, 
    1364, 
    2537, 
    1967, 
    2993, 
    2460, 
    2028, 
    1364, 
    2603, 
    2993, 
    5896, 
    5458, 
    4621, 
    1977, 
    4574, 
    848, 
    4621, 
    2028, 
    848, 
    3384, 
    4621, 
    1728, 
    1435, 
    2536, 
    5324, 
    2941, 
    2536, 
    4972, 
    5324, 
    4819, 
    4972, 
    2357, 
    5324, 
    5345, 
    5428, 
    4247, 
    5224, 
    1987, 
    770, 
    5345, 
    5093, 
    2744, 
    3111, 
    5428, 
    2744, 
    4247, 
    4455, 
    5345, 
    4455, 
    1300, 
    5245, 
    6221, 
    6504, 
    4647, 
    3797, 
    2242, 
    909, 
    143, 
    3797, 
    909, 
    1224, 
    2242, 
    3797, 
    2560, 
    1447, 
    1720, 
    2242, 
    2156, 
    1079, 
    1568, 
    1261, 
    2560, 
    2357, 
    1401, 
    603, 
    1834, 
    2357, 
    149, 
    1435, 
    6504, 
    5959, 
    1834, 
    2941, 
    5324, 
    4829, 
    6038, 
    2560, 
    4819, 
    5324, 
    2536, 
    1834, 
    1079, 
    6038, 
    4829, 
    2536, 
    2941, 
    6129, 
    1728, 
    2536, 
    4829, 
    6129, 
    2536, 
    932, 
    1728, 
    6129, 
    765, 
    6188, 
    2721, 
    5134, 
    1044, 
    967, 
    6597, 
    5134, 
    967, 
    163, 
    607, 
    5134, 
    4425, 
    1199, 
    3983, 
    1834, 
    887, 
    2242, 
    3332, 
    743, 
    2561, 
    1102, 
    1851, 
    2016, 
    2172, 
    1102, 
    1343, 
    2328, 
    2172, 
    1343, 
    1588, 
    3513, 
    3584, 
    4643, 
    715, 
    1851, 
    2172, 
    4643, 
    1102, 
    695, 
    715, 
    4643, 
    1649, 
    825, 
    2371, 
    1577, 
    5551, 
    1601, 
    3811, 
    5190, 
    2382, 
    2840, 
    1296, 
    1841, 
    1751, 
    2135, 
    4004, 
    4004, 
    1542, 
    4813, 
    4004, 
    2135, 
    1542, 
    1408, 
    4004, 
    1296, 
    1408, 
    1751, 
    4004, 
    4425, 
    162, 
    1199, 
    1044, 
    4425, 
    2135, 
    1044, 
    607, 
    4425, 
    5787, 
    632, 
    330, 
    722, 
    5787, 
    330, 
    2490, 
    6172, 
    5787, 
    3437, 
    2929, 
    2040, 
    2500, 
    3437, 
    1387, 
    734, 
    2929, 
    3437, 
    2518, 
    632, 
    5787, 
    6172, 
    2518, 
    5787, 
    3733, 
    6172, 
    2490, 
    3733, 
    1387, 
    6172, 
    875, 
    331, 
    2518, 
    5787, 
    722, 
    2490, 
    332, 
    875, 
    5223, 
    76, 
    6645, 
    77, 
    6645, 
    78, 
    77, 
    6133, 
    6645, 
    76, 
    6133, 
    79, 
    6645, 
    5030, 
    6133, 
    76, 
    74, 
    73, 
    1293, 
    1293, 
    75, 
    74, 
    1080, 
    1293, 
    73, 
    76, 
    75, 
    1293, 
    6668, 
    71, 
    70, 
    1695, 
    70, 
    594, 
    1695, 
    1080, 
    72, 
    1375, 
    1695, 
    594, 
    1375, 
    864, 
    1695, 
    69, 
    1375, 
    594, 
    6133, 
    80, 
    79, 
    78, 
    6645, 
    79, 
    5030, 
    1050, 
    6133, 
    712, 
    1953, 
    5437, 
    82, 
    4078, 
    5667, 
    1953, 
    1246, 
    5013, 
    5437, 
    1953, 
    5013, 
    1674, 
    5437, 
    1050, 
    1674, 
    712, 
    5437, 
    2509, 
    1276, 
    1975, 
    5403, 
    2446, 
    3263, 
    5403, 
    1554, 
    2446, 
    4396, 
    4936, 
    3950, 
    1582, 
    2463, 
    748, 
    5309, 
    3538, 
    3497, 
    4081, 
    5309, 
    3497, 
    3960, 
    3970, 
    5309, 
    4865, 
    4296, 
    5992, 
    4693, 
    4865, 
    3692, 
    4502, 
    4296, 
    4865, 
    3397, 
    4693, 
    3692, 
    3525, 
    3804, 
    4502, 
    3970, 
    3704, 
    5309, 
    4773, 
    3704, 
    4083, 
    3406, 
    3228, 
    3704, 
    1975, 
    2827, 
    2509, 
    748, 
    2463, 
    2827, 
    6668, 
    70, 
    1695, 
    72, 
    6668, 
    1695, 
    72, 
    71, 
    6668, 
    1080, 
    73, 
    72, 
    1674, 
    1080, 
    864, 
    712, 
    1674, 
    864, 
    5030, 
    76, 
    1293, 
    1050, 
    5030, 
    1674, 
    1050, 
    80, 
    6133, 
    1674, 
    5030, 
    1080, 
    5170, 
    1375, 
    69, 
    4596, 
    5170, 
    1733, 
    4596, 
    1554, 
    5170, 
    864, 
    1375, 
    1554, 
    864, 
    1080, 
    1695, 
    6659, 
    80, 
    6325, 
    81, 
    6659, 
    82, 
    81, 
    80, 
    6659, 
    1293, 
    1080, 
    5030, 
    3878, 
    5839, 
    6362, 
    4996, 
    5138, 
    2443, 
    3631, 
    724, 
    1564, 
    3899, 
    3631, 
    1564, 
    1797, 
    724, 
    3631, 
    1659, 
    2548, 
    4325, 
    4128, 
    4602, 
    2061, 
    4968, 
    844, 
    4325, 
    4602, 
    912, 
    2061, 
    926, 
    4602, 
    1717, 
    926, 
    2741, 
    4602, 
    4030, 
    948, 
    1190, 
    2417, 
    4030, 
    1910, 
    1921, 
    948, 
    4030, 
    6418, 
    2485, 
    5512, 
    5881, 
    2657, 
    5631, 
    5664, 
    4390, 
    4591, 
    2901, 
    5664, 
    2485, 
    5631, 
    4390, 
    5664, 
    3041, 
    3374, 
    5633, 
    5631, 
    5664, 
    2901, 
    5925, 
    6307, 
    2657, 
    5664, 
    6455, 
    2485, 
    5510, 
    4591, 
    4390, 
    6307, 
    5510, 
    4390, 
    4088, 
    3822, 
    5510, 
    2455, 
    2873, 
    5254, 
    1921, 
    3554, 
    5793, 
    5980, 
    6526, 
    2901, 
    2485, 
    6418, 
    2901, 
    5843, 
    5630, 
    6526, 
    1672, 
    6446, 
    5349, 
    6526, 
    3241, 
    2901, 
    5843, 
    6526, 
    5980, 
    5636, 
    3241, 
    6526, 
    6049, 
    3554, 
    1921, 
    1452, 
    6388, 
    1921, 
    3374, 
    3041, 
    6049, 
    5881, 
    3241, 
    3554, 
    6049, 
    5881, 
    3554, 
    3041, 
    2657, 
    5881, 
    5843, 
    2644, 
    2648, 
    5636, 
    6526, 
    5630, 
    6418, 
    5512, 
    2644, 
    5980, 
    6418, 
    5843, 
    5980, 
    2901, 
    6418, 
    2505, 
    3410, 
    3707, 
    862, 
    1278, 
    1672, 
    6119, 
    2433, 
    5572, 
    6119, 
    2853, 
    2433, 
    4264, 
    6119, 
    2599, 
    4264, 
    4471, 
    6119, 
    5534, 
    3202, 
    2853, 
    5191, 
    5534, 
    4471, 
    5191, 
    3516, 
    5534, 
    5534, 
    3516, 
    3202, 
    4562, 
    5191, 
    4471, 
    6118, 
    3516, 
    5191, 
    4830, 
    6118, 
    5191, 
    4830, 
    4917, 
    6118, 
    4054, 
    3796, 
    4917, 
    1848, 
    4054, 
    1099, 
    1848, 
    2369, 
    4278, 
    2443, 
    5138, 
    1417, 
    3680, 
    4842, 
    4996, 
    4054, 
    1848, 
    4278, 
    4487, 
    4054, 
    4278, 
    4487, 
    3796, 
    4054, 
    4663, 
    6386, 
    3516, 
    5489, 
    5946, 
    4487, 
    4278, 
    5489, 
    4487, 
    6350, 
    4671, 
    5730, 
    6379, 
    6197, 
    6318, 
    4487, 
    5946, 
    4663, 
    5489, 
    5658, 
    6197, 
    3263, 
    2446, 
    2921, 
    3497, 
    3538, 
    2921, 
    5403, 
    1953, 
    712, 
    3228, 
    3570, 
    3263, 
    3228, 
    2881, 
    3570, 
    1554, 
    1375, 
    5170, 
    864, 
    1554, 
    712, 
    5170, 
    69, 
    1733, 
    2565, 
    888, 
    2048, 
    4396, 
    3950, 
    2565, 
    1220, 
    5339, 
    2048, 
    4936, 
    1276, 
    3950, 
    2048, 
    5339, 
    4396, 
    2597, 
    1975, 
    4936, 
    2279, 
    1733, 
    2961, 
    2864, 
    2279, 
    1276, 
    3878, 
    6362, 
    1303, 
    3950, 
    2961, 
    2565, 
    5181, 
    68, 
    2294, 
    1733, 
    5181, 
    2961, 
    1733, 
    69, 
    5181, 
    2864, 
    4596, 
    2279, 
    69, 
    68, 
    5181, 
    3067, 
    2151, 
    1564, 
    2167, 
    3887, 
    3399, 
    4476, 
    4549, 
    2597, 
    3399, 
    3887, 
    2688, 
    2167, 
    1582, 
    3887, 
    5292, 
    5607, 
    6271, 
    2474, 
    5059, 
    3507, 
    6435, 
    5587, 
    5474, 
    6012, 
    6435, 
    5584, 
    6012, 
    4919, 
    6552, 
    2890, 
    4919, 
    2474, 
    6469, 
    4572, 
    5752, 
    4296, 
    4502, 
    3804, 
    3212, 
    3663, 
    3934, 
    4518, 
    3397, 
    2167, 
    4852, 
    4681, 
    4518, 
    1846, 
    4852, 
    1096, 
    3212, 
    4681, 
    4852, 
    4681, 
    4693, 
    4518, 
    4065, 
    4083, 
    4296, 
    2463, 
    3397, 
    3692, 
    2862, 
    3362, 
    3663, 
    4518, 
    2167, 
    1096, 
    4693, 
    4502, 
    4865, 
    4518, 
    4693, 
    3397, 
    4681, 
    4502, 
    4693, 
    1096, 
    4852, 
    4518, 
    3525, 
    4502, 
    4681, 
    2463, 
    1582, 
    3397, 
    1846, 
    2367, 
    2862, 
    3887, 
    4352, 
    2688, 
    4352, 
    1073, 
    2688, 
    1582, 
    4549, 
    3887, 
    1827, 
    1073, 
    4352, 
    4476, 
    1827, 
    4352, 
    4549, 
    4476, 
    4352, 
    3887, 
    4549, 
    4352, 
    1582, 
    748, 
    4549, 
    6515, 
    4936, 
    4396, 
    2597, 
    6515, 
    5525, 
    2597, 
    4936, 
    6515, 
    1975, 
    2597, 
    748, 
    1975, 
    1276, 
    4936, 
    676, 
    1534, 
    1827, 
    1534, 
    2128, 
    1073, 
    1827, 
    1534, 
    1073, 
    676, 
    3261, 
    3757, 
    2554, 
    689, 
    1541, 
    2070, 
    1429, 
    3786, 
    1230, 
    1641, 
    1940, 
    2953, 
    2554, 
    3189, 
    689, 
    2953, 
    1940, 
    2554, 
    3596, 
    3189, 
    2204, 
    1983, 
    762, 
    2246, 
    2204, 
    1230, 
    1159, 
    1983, 
    2204, 
    2177, 
    1598, 
    4093, 
    4170, 
    2830, 
    3180, 
    5108, 
    2177, 
    1112, 
    1336, 
    5108, 
    1112, 
    689, 
    816, 
    5108, 
    5727, 
    4199, 
    6173, 
    4310, 
    5727, 
    4511, 
    4411, 
    4199, 
    5727, 
    4093, 
    4609, 
    4310, 
    5686, 
    3991, 
    2833, 
    4609, 
    6532, 
    4411, 
    4217, 
    3991, 
    5686, 
    5009, 
    2877, 
    1362, 
    3352, 
    5009, 
    2336, 
    1013, 
    2877, 
    5009, 
    3034, 
    1202, 
    5143, 
    2647, 
    2425, 
    1919, 
    844, 
    2647, 
    1659, 
    844, 
    4383, 
    5697, 
    3293, 
    3597, 
    4060, 
    3867, 
    3296, 
    2749, 
    4281, 
    4060, 
    3597, 
    5867, 
    4342, 
    4668, 
    4281, 
    5867, 
    4489, 
    2749, 
    4342, 
    5867, 
    2740, 
    3991, 
    6259, 
    2833, 
    3991, 
    2740, 
    1292, 
    2288, 
    3799, 
    3293, 
    3603, 
    3597, 
    1747, 
    3293, 
    3799, 
    1747, 
    962, 
    3293, 
    3700, 
    1513, 
    2118, 
    3108, 
    3183, 
    2833, 
    3108, 
    2425, 
    3183, 
    3034, 
    2647, 
    1919, 
    1202, 
    3034, 
    1919, 
    2219, 
    1659, 
    3034, 
    3700, 
    2118, 
    2675, 
    4199, 
    2833, 
    3968, 
    1292, 
    4431, 
    1983, 
    4281, 
    3597, 
    3867, 
    6259, 
    4060, 
    4281, 
    2740, 
    6259, 
    4281, 
    4217, 
    6159, 
    6259, 
    3799, 
    3293, 
    4060, 
    5060, 
    4588, 
    2824, 
    2095, 
    5060, 
    3603, 
    2095, 
    1466, 
    5060, 
    2228, 
    4342, 
    2555, 
    1747, 
    3799, 
    2288, 
    4489, 
    2740, 
    4281, 
    3867, 
    5867, 
    4281, 
    4342, 
    1202, 
    4668, 
    2425, 
    3108, 
    1919, 
    2425, 
    1513, 
    3183, 
    1292, 
    1894, 
    2288, 
    3226, 
    4638, 
    1960, 
    2877, 
    2025, 
    1362, 
    2336, 
    5009, 
    1362, 
    2118, 
    1513, 
    4383, 
    2675, 
    2118, 
    1013, 
    1787, 
    3180, 
    1013, 
    5436, 
    3968, 
    3700, 
    2830, 
    5436, 
    2675, 
    6173, 
    4199, 
    3968, 
    4691, 
    6173, 
    5436, 
    4691, 
    4511, 
    6173, 
    4134, 
    6168, 
    2830, 
    4511, 
    5727, 
    6173, 
    5195, 
    1983, 
    4431, 
    4310, 
    4609, 
    4411, 
    762, 
    1983, 
    4609, 
    5686, 
    2833, 
    4199, 
    3108, 
    2833, 
    2740, 
    2958, 
    1112, 
    5062, 
    762, 
    4093, 
    1598, 
    4925, 
    3873, 
    2559, 
    2958, 
    4925, 
    2559, 
    4310, 
    4511, 
    4925, 
    762, 
    4609, 
    4093, 
    6168, 
    4691, 
    2830, 
    3873, 
    6168, 
    4134, 
    4511, 
    4691, 
    6168, 
    4411, 
    5727, 
    4310, 
    6173, 
    3968, 
    5436, 
    3183, 
    3968, 
    2833, 
    4925, 
    6168, 
    3873, 
    2118, 
    4383, 
    2877, 
    4638, 
    1255, 
    1960, 
    2025, 
    4638, 
    1362, 
    2025, 
    4968, 
    4638, 
    1013, 
    2118, 
    2877, 
    4968, 
    4325, 
    2265, 
    1255, 
    4968, 
    2265, 
    2025, 
    844, 
    4968, 
    1043, 
    1336, 
    1858, 
    6147, 
    2790, 
    4149, 
    4134, 
    6147, 
    4149, 
    4345, 
    4558, 
    6147, 
    2830, 
    4345, 
    4134, 
    4558, 
    3148, 
    2790, 
    4170, 
    4558, 
    4345, 
    4170, 
    2324, 
    4558, 
    1787, 
    4170, 
    3180, 
    2324, 
    1340, 
    4558, 
    816, 
    1598, 
    2177, 
    4411, 
    5686, 
    4199, 
    6532, 
    4217, 
    5686, 
    4411, 
    6532, 
    5686, 
    5195, 
    4431, 
    6532, 
    3799, 
    4431, 
    1292, 
    3799, 
    4060, 
    6159, 
    6159, 
    4060, 
    6259, 
    4431, 
    6159, 
    4217, 
    4431, 
    3799, 
    6159, 
    2988, 
    2048, 
    888, 
    1163, 
    3466, 
    3325, 
    1220, 
    2048, 
    2988, 
    3466, 
    4381, 
    1220, 
    1895, 
    2407, 
    4456, 
    1645, 
    3261, 
    4381, 
    5525, 
    1827, 
    4476, 
    2597, 
    5525, 
    4476, 
    6285, 
    1935, 
    1827, 
    5339, 
    6285, 
    5525, 
    5339, 
    1220, 
    6285, 
    6644, 
    83, 
    82, 
    1396, 
    6644, 
    82, 
    84, 
    83, 
    6644, 
    3763, 
    85, 
    84, 
    6600, 
    121, 
    120, 
    1836, 
    6600, 
    120, 
    122, 
    121, 
    6600, 
    1864, 
    118, 
    117, 
    2097, 
    5118, 
    117, 
    971, 
    120, 
    1864, 
    118, 
    1864, 
    119, 
    110, 
    109, 
    6627, 
    6642, 
    108, 
    668, 
    6627, 
    6642, 
    111, 
    6627, 
    109, 
    6642, 
    110, 
    6627, 
    111, 
    109, 
    108, 
    6642, 
    105, 
    6580, 
    106, 
    105, 
    1439, 
    4235, 
    104, 
    103, 
    6689, 
    6689, 
    6690, 
    598, 
    104, 
    6689, 
    598, 
    103, 
    6690, 
    6689, 
    6571, 
    100, 
    597, 
    6687, 
    6697, 
    597, 
    101, 
    100, 
    6571, 
    6697, 
    101, 
    6571, 
    6687, 
    597, 
    596, 
    1404, 
    6687, 
    596, 
    6697, 
    6571, 
    597, 
    102, 
    6697, 
    6687, 
    102, 
    101, 
    6697, 
    6687, 
    1404, 
    102, 
    1404, 
    596, 
    595, 
    1439, 
    2076, 
    1118, 
    102, 
    1404, 
    103, 
    595, 
    99, 
    3759, 
    3759, 
    99, 
    98, 
    2076, 
    3759, 
    935, 
    2076, 
    1404, 
    3759, 
    98, 
    97, 
    935, 
    1439, 
    1118, 
    1026, 
    6690, 
    2054, 
    105, 
    598, 
    6690, 
    105, 
    103, 
    2054, 
    6690, 
    2076, 
    935, 
    1118, 
    2054, 
    2076, 
    1439, 
    1404, 
    595, 
    3759, 
    98, 
    935, 
    3759, 
    1528, 
    95, 
    1356, 
    2054, 
    103, 
    1404, 
    2076, 
    2054, 
    1404, 
    1439, 
    105, 
    2054, 
    96, 
    95, 
    6699, 
    4246, 
    94, 
    1496, 
    2333, 
    1356, 
    998, 
    1776, 
    4446, 
    998, 
    1118, 
    1528, 
    2333, 
    95, 
    94, 
    1356, 
    1528, 
    1118, 
    935, 
    94, 
    4246, 
    1356, 
    5994, 
    2415, 
    1269, 
    1356, 
    4246, 
    998, 
    1496, 
    2415, 
    5994, 
    768, 
    1269, 
    90, 
    6009, 
    3271, 
    1299, 
    768, 
    6009, 
    1890, 
    768, 
    2520, 
    6009, 
    3875, 
    740, 
    1326, 
    998, 
    4866, 
    1776, 
    802, 
    740, 
    3875, 
    6642, 
    668, 
    111, 
    1528, 
    935, 
    97, 
    6699, 
    1528, 
    97, 
    96, 
    6699, 
    97, 
    95, 
    1528, 
    6699, 
    1356, 
    2333, 
    1528, 
    1026, 
    1118, 
    2333, 
    1026, 
    4235, 
    1439, 
    998, 
    4446, 
    2333, 
    6580, 
    107, 
    106, 
    4235, 
    6580, 
    105, 
    4235, 
    107, 
    6580, 
    108, 
    4235, 
    1026, 
    108, 
    107, 
    4235, 
    599, 
    111, 
    668, 
    93, 
    92, 
    1496, 
    92, 
    91, 
    2415, 
    2415, 
    90, 
    1269, 
    802, 
    4866, 
    5994, 
    1496, 
    92, 
    2415, 
    2520, 
    90, 
    89, 
    995, 
    6009, 
    2520, 
    1890, 
    802, 
    1269, 
    768, 
    1890, 
    1269, 
    3606, 
    1471, 
    1575, 
    2399, 
    3606, 
    740, 
    2399, 
    1471, 
    3606, 
    1299, 
    2399, 
    1890, 
    1299, 
    1471, 
    2399, 
    599, 
    1326, 
    112, 
    1496, 
    94, 
    93, 
    90, 
    2415, 
    91, 
    4866, 
    802, 
    3875, 
    4246, 
    4866, 
    998, 
    5994, 
    1269, 
    802, 
    4246, 
    5994, 
    4866, 
    4246, 
    1496, 
    5994, 
    3875, 
    1326, 
    1776, 
    668, 
    108, 
    1026, 
    1575, 
    740, 
    3606, 
    1326, 
    1575, 
    112, 
    1326, 
    740, 
    1575, 
    668, 
    1326, 
    599, 
    3875, 
    1776, 
    4866, 
    668, 
    1776, 
    1326, 
    4446, 
    1026, 
    2333, 
    668, 
    4446, 
    1776, 
    668, 
    1026, 
    4446, 
    6643, 
    600, 
    113, 
    112, 
    6643, 
    113, 
    112, 
    2273, 
    6643, 
    6643, 
    2273, 
    114, 
    6688, 
    115, 
    114, 
    2273, 
    6688, 
    114, 
    116, 
    115, 
    6688, 
    6643, 
    114, 
    600, 
    2273, 
    116, 
    6688, 
    1575, 
    2273, 
    112, 
    2097, 
    117, 
    2273, 
    5118, 
    1755, 
    971, 
    117, 
    5118, 
    1864, 
    2097, 
    1471, 
    5118, 
    116, 
    2273, 
    117, 
    1471, 
    2290, 
    5118, 
    802, 
    1890, 
    740, 
    4265, 
    1438, 
    1083, 
    1755, 
    4265, 
    1083, 
    1493, 
    1438, 
    4265, 
    3271, 
    1493, 
    1299, 
    733, 
    934, 
    2075, 
    1471, 
    2097, 
    2273, 
    2799, 
    88, 
    87, 
    2520, 
    2799, 
    1264, 
    2520, 
    89, 
    2799, 
    88, 
    2799, 
    89, 
    6009, 
    995, 
    3271, 
    90, 
    2520, 
    768, 
    1264, 
    995, 
    2520, 
    86, 
    2268, 
    87, 
    2268, 
    853, 
    2223, 
    6009, 
    1299, 
    1890, 
    733, 
    3271, 
    995, 
    733, 
    1493, 
    3271, 
    2799, 
    87, 
    1264, 
    971, 
    1083, 
    1836, 
    2075, 
    1493, 
    733, 
    119, 
    1864, 
    120, 
    2399, 
    740, 
    1890, 
    2290, 
    1755, 
    5118, 
    1493, 
    2290, 
    1299, 
    1493, 
    1755, 
    2290, 
    1471, 
    2273, 
    1575, 
    2268, 
    1264, 
    87, 
    853, 
    2268, 
    86, 
    1721, 
    1264, 
    2268, 
    2030, 
    2223, 
    853, 
    934, 
    733, 
    1721, 
    2030, 
    4248, 
    1367, 
    995, 
    1264, 
    1721, 
    3763, 
    84, 
    1309, 
    602, 
    1524, 
    123, 
    1524, 
    602, 
    741, 
    775, 
    1524, 
    741, 
    124, 
    123, 
    1524, 
    601, 
    741, 
    602, 
    1524, 
    125, 
    124, 
    122, 
    2182, 
    601, 
    775, 
    125, 
    1524, 
    4319, 
    934, 
    2223, 
    4319, 
    2075, 
    934, 
    1913, 
    4319, 
    1194, 
    1913, 
    3171, 
    4805, 
    1438, 
    1493, 
    2075, 
    4805, 
    3171, 
    2818, 
    2075, 
    4805, 
    1438, 
    4319, 
    1913, 
    4805, 
    1083, 
    971, 
    1755, 
    2075, 
    4319, 
    4805, 
    6600, 
    1836, 
    122, 
    120, 
    971, 
    1836, 
    2290, 
    1471, 
    1299, 
    4265, 
    1755, 
    1493, 
    971, 
    1864, 
    5118, 
    2182, 
    741, 
    601, 
    1836, 
    6335, 
    122, 
    6335, 
    1083, 
    2818, 
    2182, 
    3774, 
    741, 
    995, 
    1721, 
    733, 
    4856, 
    2340, 
    1803, 
    1194, 
    4105, 
    4688, 
    1194, 
    2223, 
    6296, 
    6296, 
    2030, 
    1367, 
    1194, 
    6296, 
    4105, 
    2223, 
    2030, 
    6296, 
    4105, 
    6296, 
    1367, 
    4319, 
    2223, 
    1194, 
    1721, 
    2268, 
    2223, 
    6107, 
    1309, 
    1828, 
    853, 
    3763, 
    2030, 
    853, 
    86, 
    3763, 
    2186, 
    725, 
    1961, 
    1131, 
    2186, 
    1961, 
    1803, 
    1614, 
    2186, 
    780, 
    1614, 
    1367, 
    780, 
    1565, 
    1614, 
    126, 
    125, 
    775, 
    133, 
    132, 
    2313, 
    2313, 
    131, 
    801, 
    130, 
    801, 
    131, 
    135, 
    134, 
    1630, 
    2313, 
    134, 
    133, 
    131, 
    2313, 
    132, 
    801, 
    1630, 
    2313, 
    3855, 
    1538, 
    685, 
    1793, 
    3855, 
    685, 
    1793, 
    2331, 
    4401, 
    801, 
    2331, 
    1630, 
    2835, 
    1040, 
    2132, 
    3855, 
    4401, 
    2132, 
    5571, 
    2020, 
    1505, 
    6621, 
    128, 
    127, 
    6638, 
    6621, 
    127, 
    2020, 
    6638, 
    127, 
    130, 
    129, 
    6638, 
    129, 
    128, 
    6621, 
    6638, 
    129, 
    6621, 
    2020, 
    1354, 
    130, 
    126, 
    2020, 
    127, 
    126, 
    1505, 
    2020, 
    5571, 
    1505, 
    3185, 
    2818, 
    1083, 
    1438, 
    4805, 
    2818, 
    1438, 
    1505, 
    5605, 
    2419, 
    5605, 
    775, 
    3774, 
    3171, 
    5605, 
    3774, 
    1505, 
    775, 
    5605, 
    3774, 
    6335, 
    2818, 
    85, 
    3763, 
    86, 
    6644, 
    1396, 
    84, 
    4248, 
    780, 
    1367, 
    3763, 
    4248, 
    2030, 
    889, 
    780, 
    4248, 
    2466, 
    4780, 
    2064, 
    6107, 
    1828, 
    889, 
    4248, 
    6107, 
    889, 
    4248, 
    3763, 
    6107, 
    2553, 
    1709, 
    915, 
    1396, 
    2553, 
    1828, 
    1396, 
    82, 
    5667, 
    84, 
    1396, 
    1309, 
    5013, 
    6325, 
    1050, 
    5667, 
    4078, 
    2260, 
    1709, 
    5667, 
    2260, 
    2553, 
    1396, 
    5667, 
    82, 
    6659, 
    4078, 
    5295, 
    1803, 
    1040, 
    3503, 
    5295, 
    2835, 
    3503, 
    5391, 
    5295, 
    6317, 
    3503, 
    2835, 
    4935, 
    6317, 
    2835, 
    4935, 
    5571, 
    6317, 
    5391, 
    2419, 
    4688, 
    4856, 
    1803, 
    5295, 
    5391, 
    4856, 
    5295, 
    4688, 
    4105, 
    4856, 
    1614, 
    2340, 
    1367, 
    1614, 
    1803, 
    2340, 
    1614, 
    725, 
    2186, 
    3763, 
    1309, 
    6107, 
    5013, 
    1050, 
    5437, 
    4078, 
    5013, 
    1246, 
    6325, 
    80, 
    1050, 
    4078, 
    6325, 
    5013, 
    4078, 
    6659, 
    6325, 
    2152, 
    1565, 
    780, 
    1828, 
    4780, 
    889, 
    2466, 
    5310, 
    2152, 
    2842, 
    5387, 
    2061, 
    912, 
    2842, 
    2061, 
    3663, 
    3212, 
    2862, 
    5292, 
    5192, 
    5607, 
    5387, 
    5292, 
    6271, 
    1413, 
    5387, 
    3362, 
    2842, 
    5292, 
    5387, 
    3192, 
    5192, 
    5292, 
    5192, 
    3507, 
    5059, 
    912, 
    4180, 
    2842, 
    3934, 
    3525, 
    3212, 
    6128, 
    5059, 
    6012, 
    3362, 
    5387, 
    6271, 
    3192, 
    3507, 
    5192, 
    5059, 
    2474, 
    4919, 
    3942, 
    3673, 
    3507, 
    2842, 
    4180, 
    3192, 
    5400, 
    3517, 
    5302, 
    3673, 
    5400, 
    5302, 
    2434, 
    3205, 
    5400, 
    4919, 
    2890, 
    4275, 
    3205, 
    3517, 
    5400, 
    4303, 
    4507, 
    3649, 
    6396, 
    6163, 
    6023, 
    6403, 
    6331, 
    6264, 
    6142, 
    6404, 
    6396, 
    6506, 
    6318, 
    6428, 
    6244, 
    6506, 
    6404, 
    6244, 
    6318, 
    6506, 
    5679, 
    5519, 
    6501, 
    5387, 
    1413, 
    2061, 
    3192, 
    5292, 
    2842, 
    2862, 
    2367, 
    3362, 
    2714, 
    3416, 
    1846, 
    1096, 
    3399, 
    1846, 
    724, 
    1960, 
    5490, 
    4128, 
    5791, 
    2265, 
    3416, 
    4014, 
    6277, 
    5490, 
    1960, 
    4014, 
    3416, 
    5490, 
    4014, 
    3416, 
    2714, 
    5490, 
    1797, 
    2336, 
    3226, 
    3416, 
    6277, 
    2367, 
    1630, 
    136, 
    135, 
    2313, 
    1630, 
    134, 
    801, 
    1354, 
    2331, 
    1354, 
    801, 
    130, 
    6638, 
    2020, 
    130, 
    2132, 
    1538, 
    3855, 
    4401, 
    2835, 
    2132, 
    1793, 
    4401, 
    3855, 
    2331, 
    1354, 
    4935, 
    1630, 
    2331, 
    1793, 
    4935, 
    2835, 
    4401, 
    2331, 
    4935, 
    4401, 
    1354, 
    5571, 
    4935, 
    1040, 
    1131, 
    2132, 
    1793, 
    136, 
    1630, 
    751, 
    927, 
    1538, 
    137, 
    136, 
    685, 
    138, 
    137, 
    1431, 
    1396, 
    1828, 
    1309, 
    2553, 
    915, 
    4780, 
    5667, 
    1709, 
    2553, 
    2463, 
    4081, 
    2827, 
    2921, 
    2446, 
    2864, 
    2827, 
    3497, 
    2509, 
    5403, 
    3570, 
    1953, 
    1554, 
    5403, 
    712, 
    3263, 
    3570, 
    5403, 
    3212, 
    3525, 
    4681, 
    3570, 
    1246, 
    1953, 
    4773, 
    4606, 
    3406, 
    2260, 
    1246, 
    2881, 
    1582, 
    2167, 
    3397, 
    2597, 
    4549, 
    748, 
    6078, 
    2881, 
    3228, 
    3077, 
    6078, 
    3406, 
    4772, 
    2881, 
    6078, 
    1073, 
    2151, 
    2688, 
    2434, 
    4180, 
    1706, 
    4180, 
    3942, 
    3192, 
    1706, 
    4180, 
    912, 
    2434, 
    3942, 
    4180, 
    5791, 
    4014, 
    1255, 
    2265, 
    5791, 
    1255, 
    4128, 
    6277, 
    5791, 
    1846, 
    2862, 
    4852, 
    3970, 
    4083, 
    3704, 
    3538, 
    5309, 
    3704, 
    4296, 
    3804, 
    4065, 
    5992, 
    4296, 
    4083, 
    3970, 
    5992, 
    4083, 
    3970, 
    3960, 
    5992, 
    3960, 
    3692, 
    4865, 
    3934, 
    6534, 
    3525, 
    4379, 
    3546, 
    3822, 
    3372, 
    2890, 
    2474, 
    2655, 
    3546, 
    4275, 
    2883, 
    915, 
    2701, 
    2688, 
    3067, 
    3399, 
    4014, 
    1960, 
    1255, 
    1846, 
    3416, 
    2367, 
    2714, 
    724, 
    5490, 
    4507, 
    4687, 
    3345, 
    1616, 
    3019, 
    1788, 
    4507, 
    3345, 
    3649, 
    6307, 
    5925, 
    4303, 
    4088, 
    6307, 
    4303, 
    4390, 
    2657, 
    6307, 
    6181, 
    3374, 
    1515, 
    4687, 
    5633, 
    4676, 
    6525, 
    4507, 
    5925, 
    3019, 
    5586, 
    2624, 
    5679, 
    5486, 
    5849, 
    4780, 
    2466, 
    889, 
    2553, 
    4780, 
    1828, 
    915, 
    2064, 
    4780, 
    4284, 
    2667, 
    4083, 
    2883, 
    3231, 
    3680, 
    3231, 
    2701, 
    3077, 
    2064, 
    2883, 
    2443, 
    3406, 
    6078, 
    3228, 
    4606, 
    3077, 
    3406, 
    6278, 
    4606, 
    3049, 
    3231, 
    3077, 
    4606, 
    4671, 
    6278, 
    3049, 
    5138, 
    5489, 
    4278, 
    3231, 
    6278, 
    3680, 
    6331, 
    6551, 
    5679, 
    6561, 
    5632, 
    5792, 
    6563, 
    6445, 
    6561, 
    6551, 
    6563, 
    5755, 
    6551, 
    6409, 
    6563, 
    6508, 
    6408, 
    6445, 
    6563, 
    6508, 
    6445, 
    6553, 
    6404, 
    6506, 
    6409, 
    6537, 
    6508, 
    6409, 
    6403, 
    6537, 
    6553, 
    6428, 
    6410, 
    5474, 
    5632, 
    6408, 
    6379, 
    6244, 
    6142, 
    6386, 
    6379, 
    6142, 
    5946, 
    6197, 
    6379, 
    6410, 
    6428, 
    6429, 
    6379, 
    6318, 
    6244, 
    6197, 
    5552, 
    6318, 
    5489, 
    6197, 
    5946, 
    5658, 
    6350, 
    6197, 
    4996, 
    5658, 
    5489, 
    6350, 
    5552, 
    6197, 
    4842, 
    6350, 
    5658, 
    4842, 
    4671, 
    6350, 
    5954, 
    4492, 
    4284, 
    6043, 
    5954, 
    4284, 
    4065, 
    6043, 
    4284, 
    5917, 
    5818, 
    6043, 
    5818, 
    6410, 
    6429, 
    6350, 
    5730, 
    5552, 
    4671, 
    4492, 
    5730, 
    6278, 
    4671, 
    4842, 
    3680, 
    6278, 
    4842, 
    3231, 
    4606, 
    6278, 
    5892, 
    5917, 
    6043, 
    6410, 
    5818, 
    5670, 
    5730, 
    4492, 
    5954, 
    2667, 
    4492, 
    3049, 
    5892, 
    4065, 
    3804, 
    5741, 
    5892, 
    5567, 
    6043, 
    5818, 
    5954, 
    5741, 
    5917, 
    5892, 
    5783, 
    5670, 
    5917, 
    2443, 
    2883, 
    3680, 
    2883, 
    2701, 
    3231, 
    2701, 
    1709, 
    4772, 
    1709, 
    2701, 
    915, 
    4772, 
    2260, 
    2881, 
    2701, 
    4772, 
    3077, 
    1709, 
    2260, 
    4772, 
    2466, 
    2152, 
    889, 
    1417, 
    2466, 
    2064, 
    1417, 
    5310, 
    2466, 
    4512, 
    725, 
    5442, 
    1256, 
    1961, 
    1099, 
    1256, 
    1131, 
    1961, 
    1538, 
    2132, 
    683, 
    2223, 
    934, 
    1721, 
    2340, 
    4105, 
    1367, 
    1040, 
    2835, 
    5295, 
    2419, 
    3171, 
    1913, 
    5391, 
    3503, 
    3185, 
    2419, 
    5391, 
    3185, 
    4688, 
    4856, 
    5391, 
    1194, 
    4688, 
    1913, 
    4105, 
    2340, 
    4856, 
    3774, 
    775, 
    741, 
    6335, 
    3774, 
    2182, 
    122, 
    6335, 
    2182, 
    1836, 
    1083, 
    6335, 
    3171, 
    2419, 
    5605, 
    3185, 
    1505, 
    2419, 
    1913, 
    4688, 
    2419, 
    5571, 
    1354, 
    2020, 
    3503, 
    5571, 
    3185, 
    3503, 
    6317, 
    5571, 
    126, 
    775, 
    1505, 
    2818, 
    3171, 
    3774, 
    3497, 
    2921, 
    2509, 
    4081, 
    3960, 
    5309, 
    2827, 
    4081, 
    3497, 
    2463, 
    3692, 
    4081, 
    3538, 
    3263, 
    2921, 
    3538, 
    3228, 
    3263, 
    4081, 
    3692, 
    3960, 
    3704, 
    3228, 
    3538, 
    4773, 
    3406, 
    3704, 
    3049, 
    4773, 
    2667, 
    3049, 
    4606, 
    4773, 
    3077, 
    4772, 
    6078, 
    2881, 
    1246, 
    3570, 
    2864, 
    2509, 
    2921, 
    4596, 
    2864, 
    2446, 
    1554, 
    4596, 
    2446, 
    1733, 
    2279, 
    4596, 
    1276, 
    2509, 
    2864, 
    1975, 
    748, 
    2827, 
    4078, 
    1246, 
    2260, 
    1178, 
    4233, 
    334, 
    336, 
    2243, 
    337, 
    3168, 
    339, 
    1227, 
    339, 
    338, 
    1227, 
    2543, 
    1117, 
    1863, 
    4233, 
    1178, 
    2765, 
    5223, 
    875, 
    2929, 
    334, 
    5223, 
    1178, 
    333, 
    332, 
    5223, 
    4971, 
    2573, 
    2968, 
    5950, 
    4971, 
    2968, 
    3308, 
    5950, 
    2968, 
    3521, 
    3801, 
    5950, 
    3801, 
    4062, 
    4971, 
    6224, 
    3801, 
    3521, 
    5687, 
    6224, 
    3521, 
    4160, 
    3801, 
    6224, 
    6224, 
    4374, 
    4160, 
    3209, 
    5687, 
    3521, 
    3209, 
    2683, 
    5687, 
    3000, 
    2612, 
    4160, 
    4062, 
    4817, 
    4971, 
    1144, 
    2194, 
    665, 
    4341, 
    4130, 
    3000, 
    2359, 
    3290, 
    2950, 
    1405, 
    2055, 
    4130, 
    1698, 
    3912, 
    898, 
    3290, 
    2545, 
    2950, 
    4566, 
    5687, 
    2683, 
    3912, 
    3801, 
    4160, 
    898, 
    3912, 
    2612, 
    1698, 
    2250, 
    4062, 
    5950, 
    3308, 
    3209, 
    3336, 
    3642, 
    3865, 
    1624, 
    2123, 
    1526, 
    4341, 
    2545, 
    3290, 
    4130, 
    4341, 
    3290, 
    3336, 
    3865, 
    4341, 
    38, 
    37, 
    6599, 
    6599, 
    4792, 
    592, 
    38, 
    6599, 
    592, 
    37, 
    4792, 
    6599, 
    1198, 
    4792, 
    36, 
    5103, 
    4811, 
    1826, 
    36, 
    5103, 
    1198, 
    2255, 
    31, 
    5921, 
    35, 
    2255, 
    36, 
    31, 
    2391, 
    5921, 
    4818, 
    3457, 
    2576, 
    1257, 
    4642, 
    1198, 
    5995, 
    5237, 
    4009, 
    4642, 
    5995, 
    5703, 
    1257, 
    856, 
    5995, 
    1826, 
    1257, 
    1198, 
    2770, 
    1509, 
    929, 
    5815, 
    3745, 
    4009, 
    6131, 
    5815, 
    4009, 
    2770, 
    6131, 
    4009, 
    3307, 
    5663, 
    6131, 
    5663, 
    5733, 
    5874, 
    2967, 
    5663, 
    3307, 
    2967, 
    2572, 
    5733, 
    5815, 
    5663, 
    5874, 
    4818, 
    39, 
    4792, 
    5237, 
    5995, 
    856, 
    6131, 
    5663, 
    5815, 
    3457, 
    4818, 
    5703, 
    6660, 
    51, 
    6574, 
    52, 
    6660, 
    53, 
    52, 
    51, 
    6660, 
    6575, 
    49, 
    6574, 
    50, 
    6575, 
    51, 
    50, 
    49, 
    6575, 
    6574, 
    49, 
    48, 
    2346, 
    48, 
    869, 
    53, 
    2346, 
    1382, 
    6574, 
    48, 
    2346, 
    6660, 
    6574, 
    2346, 
    51, 
    6575, 
    6574, 
    6607, 
    55, 
    54, 
    6608, 
    6607, 
    54, 
    53, 
    6648, 
    54, 
    57, 
    56, 
    6608, 
    56, 
    55, 
    6607, 
    6607, 
    6608, 
    56, 
    54, 
    6648, 
    6608, 
    6648, 
    53, 
    6583, 
    57, 
    6648, 
    6583, 
    57, 
    6608, 
    6648, 
    6583, 
    58, 
    57, 
    1382, 
    6583, 
    53, 
    1382, 
    59, 
    6583, 
    869, 
    4942, 
    2346, 
    6589, 
    48, 
    47, 
    46, 
    6589, 
    47, 
    46, 
    869, 
    6589, 
    6572, 
    43, 
    869, 
    44, 
    6572, 
    45, 
    44, 
    43, 
    6572, 
    46, 
    6572, 
    869, 
    46, 
    45, 
    6572, 
    1830, 
    43, 
    1075, 
    59, 
    1382, 
    4942, 
    48, 
    6589, 
    869, 
    2346, 
    53, 
    6660, 
    1397, 
    4942, 
    869, 
    59, 
    58, 
    6583, 
    40, 
    39, 
    6661, 
    6661, 
    39, 
    2576, 
    41, 
    6661, 
    1075, 
    41, 
    40, 
    6661, 
    42, 
    41, 
    1075, 
    42, 
    1075, 
    43, 
    1198, 
    4642, 
    4792, 
    1826, 
    1072, 
    856, 
    36, 
    2255, 
    5103, 
    4811, 
    1139, 
    3951, 
    5921, 
    2391, 
    1876, 
    5103, 
    5921, 
    4811, 
    5103, 
    2255, 
    5921, 
    3300, 
    1444, 
    2959, 
    4811, 
    5921, 
    1876, 
    31, 
    1444, 
    2391, 
    2576, 
    1075, 
    6661, 
    6131, 
    2770, 
    3614, 
    3745, 
    5995, 
    4009, 
    3457, 
    5703, 
    3745, 
    4642, 
    1257, 
    5995, 
    5237, 
    1509, 
    2770, 
    3745, 
    5703, 
    5995, 
    856, 
    1509, 
    5237, 
    5177, 
    6400, 
    1830, 
    3457, 
    6228, 
    2576, 
    5874, 
    3745, 
    5815, 
    6383, 
    929, 
    1009, 
    6383, 
    3614, 
    929, 
    2513, 
    5961, 
    2924, 
    2513, 
    6192, 
    5961, 
    3307, 
    6131, 
    3614, 
    1072, 
    2150, 
    856, 
    2150, 
    1563, 
    2614, 
    856, 
    2150, 
    1509, 
    1072, 
    4811, 
    3951, 
    6138, 
    2526, 
    2934, 
    1541, 
    6274, 
    2934, 
    3023, 
    2526, 
    6138, 
    1254, 
    3023, 
    2636, 
    2264, 
    2526, 
    3023, 
    5108, 
    1336, 
    1541, 
    1112, 
    1858, 
    1336, 
    1641, 
    1598, 
    816, 
    1940, 
    1641, 
    816, 
    1230, 
    2204, 
    1641, 
    1432, 
    1009, 
    1805, 
    2376, 
    1432, 
    1043, 
    1858, 
    2376, 
    1043, 
    3323, 
    1112, 
    2958, 
    6287, 
    4907, 
    5863, 
    2376, 
    5050, 
    2924, 
    2376, 
    1858, 
    5050, 
    3323, 
    2958, 
    3632, 
    1858, 
    3323, 
    5050, 
    1858, 
    1112, 
    3323, 
    3614, 
    5961, 
    3307, 
    6383, 
    2924, 
    5961, 
    3614, 
    6383, 
    5961, 
    1009, 
    1432, 
    6383, 
    1432, 
    2376, 
    2924, 
    4523, 
    2970, 
    819, 
    2206, 
    4950, 
    1645, 
    4327, 
    2970, 
    4523, 
    5521, 
    5850, 
    6219, 
    6219, 
    5236, 
    4640, 
    1163, 
    1895, 
    4640, 
    4113, 
    5545, 
    4327, 
    3261, 
    676, 
    1935, 
    819, 
    3261, 
    1645, 
    819, 
    3757, 
    3261, 
    2614, 
    4635, 
    929, 
    2177, 
    5108, 
    816, 
    1805, 
    1043, 
    1432, 
    4635, 
    4417, 
    1009, 
    929, 
    4635, 
    1009, 
    2614, 
    1563, 
    4635, 
    4417, 
    1959, 
    2636, 
    1009, 
    4417, 
    1805, 
    723, 
    1959, 
    4417, 
    4058, 
    790, 
    1999, 
    1959, 
    4058, 
    1254, 
    1959, 
    3977, 
    4058, 
    2636, 
    1959, 
    1254, 
    2264, 
    3023, 
    1254, 
    1043, 
    1805, 
    2636, 
    3977, 
    1620, 
    790, 
    723, 
    3977, 
    1959, 
    723, 
    1563, 
    4908, 
    633, 
    6604, 
    342, 
    341, 
    3576, 
    633, 
    6625, 
    344, 
    343, 
    1151, 
    6625, 
    343, 
    634, 
    344, 
    6625, 
    1151, 
    345, 
    6625, 
    6625, 
    345, 
    634, 
    6175, 
    2814, 
    1410, 
    3850, 
    6175, 
    1151, 
    3850, 
    4116, 
    6175, 
    1437, 
    3576, 
    341, 
    1437, 
    933, 
    5385, 
    6665, 
    346, 
    1410, 
    347, 
    6665, 
    348, 
    347, 
    346, 
    6665, 
    6601, 
    349, 
    348, 
    350, 
    635, 
    1074, 
    6601, 
    635, 
    349, 
    1074, 
    6601, 
    348, 
    1074, 
    635, 
    6601, 
    5443, 
    1410, 
    2364, 
    2197, 
    5905, 
    1149, 
    5905, 
    348, 
    6665, 
    1149, 
    5905, 
    5443, 
    1074, 
    348, 
    5905, 
    351, 
    350, 
    1074, 
    1843, 
    2364, 
    2814, 
    6650, 
    24, 
    1377, 
    25, 
    6650, 
    591, 
    25, 
    24, 
    6650, 
    1031, 
    1377, 
    24, 
    21, 
    6663, 
    22, 
    6663, 
    590, 
    22, 
    20, 
    6664, 
    21, 
    21, 
    6664, 
    6663, 
    6674, 
    20, 
    6613, 
    6664, 
    6674, 
    23, 
    6664, 
    20, 
    6674, 
    590, 
    6664, 
    23, 
    590, 
    6663, 
    6664, 
    6613, 
    20, 
    19, 
    1031, 
    6613, 
    19, 
    23, 
    6674, 
    6613, 
    1031, 
    24, 
    6613, 
    1031, 
    19, 
    18, 
    1377, 
    1281, 
    6650, 
    4581, 
    1377, 
    18, 
    17, 
    4814, 
    18, 
    940, 
    3819, 
    4581, 
    3819, 
    2080, 
    1281, 
    4581, 
    3819, 
    1377, 
    940, 
    2080, 
    3819, 
    24, 
    23, 
    6613, 
    591, 
    6650, 
    1281, 
    6631, 
    28, 
    27, 
    6631, 
    29, 
    28, 
    6620, 
    6631, 
    27, 
    6620, 
    30, 
    6631, 
    6588, 
    26, 
    1444, 
    30, 
    6588, 
    31, 
    6587, 
    26, 
    6588, 
    6620, 
    6587, 
    30, 
    29, 
    6631, 
    30, 
    27, 
    6587, 
    6620, 
    27, 
    26, 
    6587, 
    6588, 
    30, 
    6587, 
    3977, 
    790, 
    4058, 
    4908, 
    2190, 
    3977, 
    723, 
    4908, 
    3977, 
    1563, 
    2150, 
    4908, 
    2272, 
    2734, 
    1725, 
    4811, 
    1876, 
    1139, 
    1826, 
    4811, 
    1072, 
    1826, 
    1198, 
    5103, 
    2639, 
    3877, 
    3433, 
    3977, 
    2190, 
    1620, 
    1139, 
    1876, 
    3025, 
    4814, 
    4307, 
    5548, 
    18, 
    4814, 
    4581, 
    17, 
    1185, 
    4814, 
    4740, 
    3174, 
    1970, 
    1725, 
    2734, 
    3877, 
    1268, 
    3493, 
    2272, 
    5132, 
    5071, 
    2652, 
    4634, 
    5132, 
    4990, 
    5248, 
    4236, 
    5142, 
    4589, 
    5073, 
    4761, 
    5132, 
    2652, 
    4990, 
    6360, 
    5813, 
    5661, 
    5073, 
    6360, 
    4933, 
    5073, 
    6341, 
    6361, 
    5401, 
    2652, 
    5071, 
    2639, 
    3433, 
    3723, 
    3493, 
    3777, 
    2734, 
    2272, 
    3493, 
    2734, 
    5577, 
    2822, 
    5541, 
    2639, 
    3723, 
    3025, 
    3777, 
    4991, 
    3104, 
    2734, 
    3777, 
    3104, 
    5854, 
    6248, 
    4161, 
    3914, 
    5854, 
    4161, 
    5712, 
    5558, 
    6320, 
    4389, 
    2632, 
    1317, 
    4934, 
    5073, 
    4589, 
    5431, 
    5347, 
    5968, 
    790, 
    5431, 
    4763, 
    1620, 
    4214, 
    5431, 
    5746, 
    6555, 
    6439, 
    5734, 
    5661, 
    6454, 
    5530, 
    5734, 
    5558, 
    5401, 
    5661, 
    5734, 
    5133, 
    4991, 
    5614, 
    5625, 
    5133, 
    5614, 
    4934, 
    5968, 
    6341, 
    6444, 
    4473, 
    5625, 
    4473, 
    3723, 
    5133, 
    2564, 
    4473, 
    4214, 
    5133, 
    3433, 
    4991, 
    5827, 
    6005, 
    4933, 
    4008, 
    5142, 
    4236, 
    5868, 
    4761, 
    6005, 
    4998, 
    5868, 
    5142, 
    4998, 
    4589, 
    5868, 
    2190, 
    1139, 
    2564, 
    5548, 
    4307, 
    1725, 
    940, 
    5548, 
    1725, 
    4581, 
    4814, 
    5548, 
    3174, 
    3493, 
    1268, 
    1970, 
    3174, 
    1268, 
    5746, 
    5577, 
    6555, 
    3174, 
    5577, 
    3493, 
    3174, 
    2822, 
    5577, 
    4307, 
    3922, 
    2272, 
    940, 
    4581, 
    5548, 
    4509, 
    1051, 
    3922, 
    4814, 
    4509, 
    4307, 
    1185, 
    1051, 
    4509, 
    4380, 
    2140, 
    1498, 
    1725, 
    4307, 
    2272, 
    1051, 
    2140, 
    3922, 
    3163, 
    2809, 
    5057, 
    1508, 
    3163, 
    2421, 
    3002, 
    3338, 
    3163, 
    2114, 
    3002, 
    1508, 
    3338, 
    2809, 
    3163, 
    3200, 
    5624, 
    3002, 
    6322, 
    2851, 
    2431, 
    5566, 
    6322, 
    5701, 
    5624, 
    2851, 
    6322, 
    3200, 
    2851, 
    5624, 
    1008, 
    3200, 
    2114, 
    4178, 
    1784, 
    3795, 
    5701, 
    2855, 
    5530, 
    5712, 
    5701, 
    5530, 
    5566, 
    5624, 
    6322, 
    3922, 
    1268, 
    2272, 
    4859, 
    5157, 
    1051, 
    4380, 
    1268, 
    3922, 
    2140, 
    4380, 
    3922, 
    1498, 
    699, 
    5926, 
    2202, 
    3, 
    2, 
    1, 
    2202, 
    2, 
    1, 
    1181, 
    2202, 
    6576, 
    584, 
    583, 
    582, 
    6576, 
    583, 
    582, 
    4118, 
    6576, 
    4118, 
    584, 
    6576, 
    579, 
    578, 
    1829, 
    662, 
    1829, 
    578, 
    705, 
    662, 
    577, 
    580, 
    1748, 
    581, 
    1829, 
    580, 
    579, 
    705, 
    1829, 
    662, 
    705, 
    580, 
    1829, 
    1347, 
    576, 
    575, 
    1407, 
    1631, 
    575, 
    942, 
    963, 
    1347, 
    580, 
    705, 
    1748, 
    577, 
    576, 
    963, 
    1748, 
    963, 
    1522, 
    1631, 
    942, 
    1347, 
    1126, 
    1270, 
    1021, 
    4118, 
    585, 
    584, 
    4118, 
    1522, 
    1021, 
    581, 
    1748, 
    582, 
    705, 
    963, 
    1748, 
    2499, 
    4320, 
    903, 
    5412, 
    5604, 
    2499, 
    1727, 
    942, 
    2109, 
    4320, 
    942, 
    804, 
    903, 
    4320, 
    804, 
    2109, 
    942, 
    4320, 
    1021, 
    1727, 
    1126, 
    1522, 
    942, 
    1727, 
    4118, 
    1748, 
    1522, 
    585, 
    4118, 
    1021, 
    582, 
    1748, 
    4118, 
    963, 
    942, 
    1522, 
    577, 
    963, 
    705, 
    576, 
    1347, 
    963, 
    2499, 
    903, 
    3029, 
    4679, 
    4850, 
    5412, 
    2109, 
    4320, 
    2499, 
    574, 
    1407, 
    575, 
    4293, 
    5048, 
    6024, 
    6021, 
    4293, 
    1498, 
    2140, 
    6021, 
    1498, 
    2140, 
    5157, 
    6021, 
    5180, 
    4358, 
    1000, 
    4077, 
    5048, 
    4293, 
    5399, 
    1361, 
    1853, 
    6394, 
    6222, 
    5399, 
    5280, 
    6394, 
    5301, 
    6110, 
    6222, 
    6394, 
    6222, 
    1361, 
    5399, 
    1270, 
    585, 
    1021, 
    2643, 
    2621, 
    1089, 
    3475, 
    2643, 
    1839, 
    1407, 
    3475, 
    1839, 
    5702, 
    1369, 
    5252, 
    5137, 
    3008, 
    2643, 
    1237, 
    2252, 
    1574, 
    3029, 
    1089, 
    2161, 
    2252, 
    3029, 
    2161, 
    1328, 
    2499, 
    3029, 
    1727, 
    1021, 
    1522, 
    2109, 
    1126, 
    1727, 
    1089, 
    3029, 
    903, 
    1237, 
    1000, 
    4358, 
    4928, 
    1, 
    663, 
    4928, 
    1181, 
    1, 
    2413, 
    1905, 
    4928, 
    2109, 
    2499, 
    5604, 
    4679, 
    2252, 
    1237, 
    4554, 
    4679, 
    4358, 
    1328, 
    2252, 
    4679, 
    4358, 
    4679, 
    1237, 
    6222, 
    5048, 
    4077, 
    1361, 
    6222, 
    4077, 
    5399, 
    5301, 
    6394, 
    2202, 
    5301, 
    3, 
    6394, 
    5377, 
    6110, 
    1905, 
    5280, 
    1181, 
    4554, 
    4358, 
    5377, 
    663, 
    586, 
    4928, 
    5725, 
    843, 
    2024, 
    6021, 
    5157, 
    5725, 
    4859, 
    1658, 
    5157, 
    2218, 
    1658, 
    4859, 
    17, 
    2218, 
    1185, 
    16, 
    15, 
    3366, 
    3366, 
    2069, 
    1658, 
    9, 
    6617, 
    10, 
    6617, 
    11, 
    10, 
    8, 
    6617, 
    9, 
    8, 
    6618, 
    6617, 
    6618, 
    11, 
    6617, 
    6581, 
    6618, 
    8, 
    6581, 
    11, 
    6618, 
    7, 
    6582, 
    8, 
    12, 
    11, 
    6581, 
    6582, 
    12, 
    6581, 
    8, 
    6582, 
    6581, 
    7, 
    6, 
    6582, 
    6632, 
    6, 
    6633, 
    6582, 
    6632, 
    12, 
    6582, 
    6, 
    6632, 
    6633, 
    12, 
    6632, 
    6677, 
    14, 
    13, 
    6678, 
    6677, 
    13, 
    589, 
    14, 
    6677, 
    6677, 
    6678, 
    589, 
    6633, 
    13, 
    12, 
    2069, 
    6633, 
    6, 
    2069, 
    6678, 
    6633, 
    588, 
    803, 
    4, 
    803, 
    5, 
    4, 
    803, 
    6, 
    5, 
    587, 
    1853, 
    1592, 
    5399, 
    3, 
    5301, 
    1592, 
    1853, 
    1361, 
    587, 
    3, 
    1853, 
    6024, 
    5048, 
    5180, 
    1425, 
    1361, 
    2024, 
    2069, 
    1425, 
    843, 
    1658, 
    2069, 
    843, 
    6678, 
    13, 
    6633, 
    15, 
    6678, 
    2069, 
    15, 
    589, 
    6678, 
    803, 
    1592, 
    1425, 
    5301, 
    1181, 
    5280, 
    5926, 
    699, 
    5388, 
    5725, 
    4077, 
    4293, 
    6021, 
    5725, 
    4293, 
    5157, 
    843, 
    5725, 
    3, 
    5399, 
    1853, 
    2140, 
    1051, 
    5157, 
    2024, 
    1361, 
    4077, 
    5725, 
    2024, 
    4077, 
    843, 
    1425, 
    2024, 
    6, 
    1425, 
    2069, 
    1592, 
    588, 
    587, 
    1425, 
    1592, 
    1361, 
    803, 
    588, 
    1592, 
    6, 
    803, 
    1425, 
    1181, 
    5301, 
    2202, 
    3366, 
    1658, 
    2218, 
    16, 
    3366, 
    2218, 
    15, 
    2069, 
    3366, 
    2225, 
    5252, 
    1369, 
    903, 
    1839, 
    1089, 
    1407, 
    574, 
    3475, 
    1631, 
    1407, 
    1839, 
    942, 
    1631, 
    804, 
    1347, 
    575, 
    1631, 
    574, 
    855, 
    3475, 
    2134, 
    1915, 
    1042, 
    3930, 
    2134, 
    1042, 
    4578, 
    3930, 
    1042, 
    1608, 
    5415, 
    3930, 
    1540, 
    1508, 
    2421, 
    4990, 
    2652, 
    2432, 
    4634, 
    4990, 
    2653, 
    4634, 
    4447, 
    5132, 
    2965, 
    4447, 
    3306, 
    5142, 
    4008, 
    4998, 
    2570, 
    4236, 
    4447, 
    4589, 
    2632, 
    4389, 
    4617, 
    5112, 
    2570, 
    4998, 
    2632, 
    4589, 
    4761, 
    5868, 
    4589, 
    4008, 
    3743, 
    4998, 
    3738, 
    1574, 
    2816, 
    5920, 
    2852, 
    5740, 
    2435, 
    5920, 
    5740, 
    2855, 
    2431, 
    5920, 
    3643, 
    5982, 
    3914, 
    4892, 
    6037, 
    2759, 
    5701, 
    2431, 
    2855, 
    5712, 
    5982, 
    5701, 
    3643, 
    3338, 
    5566, 
    2809, 
    3338, 
    3643, 
    2431, 
    3670, 
    5920, 
    1445, 
    2682, 
    2081, 
    1124, 
    4578, 
    4655, 
    5137, 
    2502, 
    3008, 
    3475, 
    5137, 
    2643, 
    5702, 
    855, 
    1369, 
    5137, 
    5702, 
    5252, 
    3475, 
    855, 
    5702, 
    1608, 
    773, 
    5415, 
    5252, 
    2502, 
    5137, 
    3475, 
    5702, 
    5137, 
    2225, 
    2914, 
    5252, 
    4690, 
    4655, 
    2225, 
    2682, 
    4690, 
    1369, 
    2384, 
    1867, 
    4690, 
    1197, 
    2914, 
    2225, 
    5388, 
    1000, 
    4003, 
    903, 
    804, 
    1839, 
    574, 
    2081, 
    855, 
    1631, 
    1839, 
    804, 
    1839, 
    2643, 
    1089, 
    6037, 
    5039, 
    2809, 
    1197, 
    3917, 
    2914, 
    5057, 
    2809, 
    5039, 
    3917, 
    5057, 
    5039, 
    1915, 
    2421, 
    5057, 
    5057, 
    2421, 
    3163, 
    2621, 
    2816, 
    2161, 
    1089, 
    2621, 
    2161, 
    5401, 
    2435, 
    5740, 
    4933, 
    6360, 
    5071, 
    6424, 
    2822, 
    4567, 
    6424, 
    5541, 
    2822, 
    6248, 
    6424, 
    4375, 
    6248, 
    6313, 
    6424, 
    4161, 
    6248, 
    4375, 
    5854, 
    5712, 
    6320, 
    2435, 
    5734, 
    5530, 
    5948, 
    5813, 
    6361, 
    6439, 
    4991, 
    3777, 
    5746, 
    6439, 
    3777, 
    6425, 
    5614, 
    6439, 
    4740, 
    2822, 
    3174, 
    739, 
    4740, 
    1970, 
    739, 
    3738, 
    4740, 
    5566, 
    5982, 
    3643, 
    6313, 
    6320, 
    6236, 
    5982, 
    5712, 
    5854, 
    3914, 
    5982, 
    5854, 
    5566, 
    5701, 
    5982, 
    5530, 
    5558, 
    5712, 
    5401, 
    5734, 
    2435, 
    6381, 
    5813, 
    5948, 
    6545, 
    6236, 
    6454, 
    5813, 
    6545, 
    6454, 
    6381, 
    6438, 
    6545, 
    5614, 
    6381, 
    5948, 
    6438, 
    6313, 
    6545, 
    6424, 
    6313, 
    5541, 
    6320, 
    5558, 
    6236, 
    6248, 
    6320, 
    6313, 
    6248, 
    5854, 
    6320, 
    5558, 
    5734, 
    6454, 
    4567, 
    4375, 
    6424, 
    4740, 
    4567, 
    2822, 
    3738, 
    3450, 
    4567, 
    3450, 
    3124, 
    4375, 
    3124, 
    2759, 
    4161, 
    5462, 
    4571, 
    3124, 
    2643, 
    3008, 
    2621, 
    2502, 
    4378, 
    4571, 
    3917, 
    1197, 
    1915, 
    4378, 
    2914, 
    3917, 
    5039, 
    4892, 
    4378, 
    1915, 
    5057, 
    3917, 
    2809, 
    3643, 
    6037, 
    4571, 
    3008, 
    2502, 
    4892, 
    4571, 
    4378, 
    2759, 
    3124, 
    4571, 
    2502, 
    5252, 
    2914, 
    1042, 
    1915, 
    1197, 
    5624, 
    3338, 
    3002, 
    2431, 
    5701, 
    6322, 
    5566, 
    3338, 
    5624, 
    2435, 
    5530, 
    2855, 
    5039, 
    4378, 
    3917, 
    6037, 
    4892, 
    5039, 
    3914, 
    6037, 
    3643, 
    3914, 
    2759, 
    6037, 
    2759, 
    4571, 
    4892, 
    2502, 
    2914, 
    4378, 
    3163, 
    1508, 
    3002, 
    4003, 
    1237, 
    1574, 
    739, 
    4003, 
    1574, 
    739, 
    5388, 
    4003, 
    5180, 
    1000, 
    699, 
    6024, 
    5180, 
    699, 
    1498, 
    6024, 
    699, 
    1498, 
    4293, 
    6024, 
    6110, 
    5377, 
    4358, 
    5048, 
    6110, 
    5180, 
    5048, 
    6222, 
    6110, 
    6110, 
    4358, 
    5180, 
    6394, 
    5280, 
    5377, 
    5280, 
    4554, 
    5377, 
    1905, 
    4554, 
    5280, 
    1905, 
    2413, 
    4850, 
    5604, 
    4850, 
    2413, 
    1328, 
    5412, 
    2499, 
    1328, 
    4679, 
    5412, 
    5604, 
    2413, 
    1126, 
    2109, 
    5604, 
    1126, 
    5412, 
    4850, 
    5604, 
    4554, 
    4850, 
    4679, 
    4554, 
    1905, 
    4850, 
    3029, 
    2252, 
    1328, 
    2161, 
    1574, 
    2252, 
    4003, 
    1000, 
    1237, 
    1444, 
    26, 
    1281, 
    1270, 
    1126, 
    2413, 
    4928, 
    1270, 
    2413, 
    1181, 
    4928, 
    1905, 
    586, 
    1270, 
    4928, 
    586, 
    585, 
    1270, 
    704, 
    1056, 
    5086, 
    5086, 
    370, 
    369, 
    3599, 
    5086, 
    369, 
    1056, 
    371, 
    5086, 
    3599, 
    367, 
    812, 
    3599, 
    812, 
    704, 
    368, 
    3599, 
    369, 
    368, 
    367, 
    3599, 
    640, 
    1241, 
    367, 
    2719, 
    1842, 
    1092, 
    3669, 
    3368, 
    3524, 
    3803, 
    3669, 
    3524, 
    2163, 
    1578, 
    3669, 
    5214, 
    5958, 
    2363, 
    3368, 
    3036, 
    3211, 
    3094, 
    3524, 
    3211, 
    3669, 
    1578, 
    3531, 
    6010, 
    5764, 
    3144, 
    6309, 
    6010, 
    5524, 
    5600, 
    5764, 
    6010, 
    5308, 
    3227, 
    4055, 
    2058, 
    5308, 
    908, 
    2880, 
    3227, 
    5308, 
    5958, 
    2880, 
    1409, 
    2363, 
    5958, 
    1409, 
    5214, 
    2785, 
    6471, 
    3227, 
    2462, 
    4055, 
    5958, 
    6471, 
    2880, 
    6010, 
    3144, 
    2685, 
    6471, 
    5764, 
    5600, 
    2880, 
    6471, 
    5600, 
    5958, 
    5214, 
    6471, 
    2785, 
    3144, 
    5764, 
    4018, 
    3396, 
    3065, 
    4209, 
    4018, 
    5494, 
    2650, 
    4767, 
    2442, 
    1148, 
    4018, 
    4209, 
    1148, 
    890, 
    4018, 
    4407, 
    812, 
    1241, 
    2462, 
    5876, 
    1241, 
    4191, 
    704, 
    4407, 
    5876, 
    3227, 
    5600, 
    3959, 
    2625, 
    4191, 
    1409, 
    703, 
    4851, 
    4055, 
    364, 
    908, 
    5360, 
    800, 
    5155, 
    372, 
    2005, 
    681, 
    372, 
    1056, 
    2005, 
    571, 
    2081, 
    572, 
    2081, 
    571, 
    1445, 
    573, 
    2081, 
    574, 
    573, 
    572, 
    2081, 
    6702, 
    470, 
    469, 
    649, 
    6590, 
    469, 
    6702, 
    471, 
    470, 
    6590, 
    6702, 
    469, 
    6590, 
    471, 
    6702, 
    6591, 
    6590, 
    649, 
    468, 
    6591, 
    649, 
    472, 
    6590, 
    6591, 
    472, 
    471, 
    6590, 
    6591, 
    468, 
    6614, 
    6614, 
    472, 
    6591, 
    6615, 
    6614, 
    468, 
    6615, 
    472, 
    6614, 
    6615, 
    473, 
    472, 
    467, 
    6615, 
    468, 
    6673, 
    6120, 
    473, 
    467, 
    6673, 
    6615, 
    467, 
    6120, 
    6673, 
    2372, 
    3895, 
    4519, 
    2099, 
    975, 
    4844, 
    4695, 
    1760, 
    2587, 
    2274, 
    1726, 
    975, 
    6693, 
    2274, 
    464, 
    463, 
    6693, 
    464, 
    6616, 
    459, 
    6693, 
    459, 
    458, 
    2274, 
    5666, 
    1305, 
    1446, 
    5422, 
    4695, 
    2587, 
    5422, 
    4868, 
    4695, 
    3766, 
    5422, 
    2587, 
    4977, 
    4868, 
    5422, 
    3480, 
    4977, 
    3766, 
    3480, 
    2089, 
    4977, 
    952, 
    1739, 
    4868, 
    2296, 
    1305, 
    4033, 
    941, 
    2296, 
    1760, 
    941, 
    2082, 
    2296, 
    4001, 
    4227, 
    5165, 
    2748, 
    3115, 
    3415, 
    1712, 
    2262, 
    3089, 
    2574, 
    3294, 
    3598, 
    5528, 
    5743, 
    3588, 
    1589, 
    1070, 
    474, 
    6120, 
    5207, 
    2173, 
    6615, 
    6673, 
    473, 
    467, 
    5080, 
    6120, 
    4022, 
    3246, 
    3557, 
    2283, 
    3088, 
    1283, 
    3895, 
    1852, 
    3088, 
    4519, 
    1421, 
    2372, 
    1739, 
    4519, 
    3895, 
    952, 
    2089, 
    4774, 
    1421, 
    5414, 
    3604, 
    3995, 
    2524, 
    2501, 
    6074, 
    4133, 
    4223, 
    3297, 
    3604, 
    3995, 
    1852, 
    3297, 
    3122, 
    3604, 
    2524, 
    3995, 
    2372, 
    3604, 
    3297, 
    2372, 
    1421, 
    3604, 
    4774, 
    2066, 
    1421, 
    4519, 
    4774, 
    1421, 
    2089, 
    1456, 
    5653, 
    2904, 
    5882, 
    2489, 
    5565, 
    4119, 
    6169, 
    6430, 
    4329, 
    5565, 
    923, 
    1690, 
    4329, 
    4213, 
    3245, 
    3556, 
    5478, 
    4213, 
    3987, 
    6436, 
    2535, 
    5882, 
    4427, 
    6436, 
    5882, 
    5585, 
    3232, 
    6436, 
    4519, 
    952, 
    4774, 
    3089, 
    3115, 
    1712, 
    3711, 
    2748, 
    3415, 
    3103, 
    3711, 
    2733, 
    3103, 
    3432, 
    3976, 
    5414, 
    1421, 
    2066, 
    3256, 
    5414, 
    3564, 
    3256, 
    2524, 
    5414, 
    3711, 
    3976, 
    5596, 
    2524, 
    3604, 
    5414, 
    2173, 
    3246, 
    4022, 
    4022, 
    3557, 
    3830, 
    1589, 
    4022, 
    1070, 
    1589, 
    2173, 
    4022, 
    1103, 
    3246, 
    2173, 
    4022, 
    1561, 
    1070, 
    2755, 
    3557, 
    3246, 
    2755, 
    2556, 
    6282, 
    2905, 
    779, 
    1992, 
    5207, 
    5080, 
    3088, 
    1589, 
    6120, 
    2173, 
    6120, 
    5080, 
    5207, 
    465, 
    1475, 
    466, 
    3088, 
    1852, 
    1103, 
    2173, 
    5207, 
    1103, 
    2283, 
    1739, 
    3895, 
    2099, 
    4844, 
    1283, 
    3895, 
    2372, 
    1852, 
    2283, 
    3895, 
    3088, 
    1739, 
    952, 
    4519, 
    6267, 
    975, 
    4695, 
    2283, 
    4844, 
    6267, 
    2283, 
    1283, 
    4844, 
    465, 
    2099, 
    1475, 
    464, 
    2274, 
    2099, 
    6679, 
    447, 
    446, 
    1215, 
    6679, 
    446, 
    448, 
    447, 
    6679, 
    455, 
    3839, 
    456, 
    647, 
    679, 
    451, 
    679, 
    452, 
    451, 
    955, 
    854, 
    4793, 
    450, 
    955, 
    647, 
    450, 
    449, 
    1506, 
    453, 
    452, 
    679, 
    454, 
    453, 
    1459, 
    4793, 
    1459, 
    453, 
    955, 
    4793, 
    679, 
    854, 
    1459, 
    4793, 
    2087, 
    1665, 
    950, 
    710, 
    2087, 
    874, 
    1454, 
    1195, 
    2087, 
    456, 
    3839, 
    648, 
    2087, 
    950, 
    874, 
    647, 
    955, 
    679, 
    4459, 
    449, 
    448, 
    2303, 
    4459, 
    1215, 
    1506, 
    449, 
    4459, 
    854, 
    1506, 
    950, 
    955, 
    450, 
    1506, 
    1665, 
    854, 
    950, 
    3839, 
    1665, 
    1195, 
    648, 
    3839, 
    1195, 
    455, 
    1459, 
    3839, 
    1459, 
    854, 
    1665, 
    454, 
    1459, 
    455, 
    453, 
    679, 
    4793, 
    3064, 
    950, 
    1506, 
    4459, 
    3064, 
    1506, 
    2303, 
    1682, 
    3064, 
    1446, 
    1682, 
    1061, 
    874, 
    950, 
    1682, 
    3839, 
    1459, 
    1665, 
    1125, 
    1215, 
    446, 
    1446, 
    1061, 
    774, 
    2303, 
    3064, 
    4459, 
    1061, 
    2303, 
    1215, 
    1061, 
    1682, 
    2303, 
    1125, 
    1609, 
    1215, 
    1454, 
    648, 
    1195, 
    1125, 
    446, 
    445, 
    753, 
    5141, 
    445, 
    1609, 
    1061, 
    1215, 
    461, 
    460, 
    6567, 
    6567, 
    460, 
    6566, 
    462, 
    6567, 
    6566, 
    462, 
    461, 
    6567, 
    6616, 
    460, 
    459, 
    6616, 
    6566, 
    460, 
    2274, 
    6693, 
    459, 
    463, 
    6566, 
    6616, 
    463, 
    462, 
    6566, 
    6693, 
    463, 
    6616, 
    1726, 
    941, 
    1760, 
    2099, 
    2274, 
    975, 
    458, 
    1386, 
    1726, 
    1386, 
    458, 
    457, 
    648, 
    1454, 
    457, 
    710, 
    941, 
    1386, 
    1454, 
    710, 
    1386, 
    457, 
    1454, 
    1386, 
    1195, 
    1665, 
    2087, 
    1454, 
    2087, 
    710, 
    955, 
    1506, 
    854, 
    1215, 
    448, 
    6679, 
    1682, 
    950, 
    3064, 
    4459, 
    448, 
    1215, 
    1446, 
    1305, 
    2082, 
    1682, 
    1446, 
    874, 
    6456, 
    3129, 
    2766, 
    4033, 
    6456, 
    5671, 
    5666, 
    3129, 
    6456, 
    774, 
    5666, 
    1446, 
    774, 
    3129, 
    5666, 
    1609, 
    774, 
    1061, 
    5713, 
    3808, 
    4070, 
    5803, 
    5713, 
    4070, 
    5141, 
    753, 
    5713, 
    445, 
    5141, 
    1125, 
    753, 
    3808, 
    5713, 
    6148, 
    1587, 
    1172, 
    4070, 
    3808, 
    6148, 
    6541, 
    4070, 
    2649, 
    6541, 
    6449, 
    5803, 
    3035, 
    6541, 
    2649, 
    5674, 
    6449, 
    6541, 
    5652, 
    6448, 
    5803, 
    3035, 
    5674, 
    6541, 
    2449, 
    5304, 
    6448, 
    6164, 
    5304, 
    1609, 
    5713, 
    6164, 
    5141, 
    6448, 
    5304, 
    6164, 
    753, 
    1587, 
    3808, 
    5653, 
    3838, 
    2066, 
    4774, 
    5653, 
    2066, 
    4774, 
    2089, 
    5653, 
    5653, 
    1456, 
    3838, 
    1760, 
    2296, 
    2587, 
    5996, 
    2766, 
    5042, 
    2089, 
    952, 
    4977, 
    2587, 
    2296, 
    4033, 
    3838, 
    4536, 
    918, 
    6148, 
    3808, 
    1587, 
    1101, 
    6148, 
    1172, 
    2903, 
    3244, 
    6253, 
    5042, 
    2867, 
    4895, 
    6385, 
    5996, 
    5042, 
    4825, 
    6385, 
    4895, 
    4825, 
    3480, 
    6385, 
    2766, 
    2449, 
    5042, 
    6164, 
    1125, 
    5141, 
    5585, 
    4213, 
    5478, 
    2535, 
    6436, 
    3232, 
    4427, 
    4213, 
    5585, 
    6436, 
    4427, 
    5585, 
    2467, 
    6039, 
    2535, 
    2904, 
    4427, 
    5882, 
    3245, 
    4213, 
    4427, 
    6169, 
    3853, 
    6052, 
    5565, 
    4329, 
    4119, 
    2489, 
    5565, 
    2904, 
    6430, 
    5569, 
    923, 
    2489, 
    6430, 
    5565, 
    2489, 
    5569, 
    6430, 
    6075, 
    885, 
    1253, 
    4329, 
    6075, 
    4119, 
    4329, 
    1690, 
    6075, 
    5098, 
    3432, 
    4958, 
    5478, 
    3722, 
    5098, 
    3541, 
    5585, 
    5478, 
    3556, 
    3829, 
    3987, 
    4205, 
    4095, 
    5366, 
    3829, 
    4095, 
    3722, 
    3829, 
    5169, 
    4095, 
    3987, 
    3829, 
    3722, 
    3829, 
    6052, 
    5169, 
    6052, 
    3581, 
    5169, 
    3245, 
    6052, 
    3556, 
    3853, 
    3581, 
    6052, 
    2904, 
    5565, 
    6169, 
    5816, 
    1253, 
    4711, 
    4205, 
    3976, 
    3432, 
    3722, 
    4205, 
    3432, 
    4095, 
    2501, 
    5366, 
    2550, 
    5618, 
    2955, 
    3616, 
    6434, 
    2550, 
    5780, 
    5914, 
    5721, 
    5505, 
    5780, 
    5721, 
    6460, 
    5509, 
    5695, 
    6461, 
    6460, 
    6365, 
    6544, 
    5509, 
    6460, 
    5492, 
    5999, 
    3988, 
    5682, 
    5644, 
    5492, 
    6200, 
    5914, 
    6040, 
    4804, 
    3435, 
    3106, 
    4958, 
    4804, 
    3106, 
    3103, 
    2733, 
    4804, 
    5028, 
    3415, 
    3089, 
    5165, 
    5028, 
    3089, 
    4441, 
    2733, 
    5028, 
    2574, 
    2969, 
    3294, 
    4964, 
    6474, 
    2591, 
    6457, 
    5676, 
    6411, 
    4723, 
    6457, 
    5735, 
    4636, 
    5676, 
    6457, 
    5602, 
    3573, 
    5470, 
    5172, 
    4035, 
    1065, 
    3114, 
    5036, 
    3443, 
    3868, 
    4131, 
    4259, 
    2956, 
    5693, 
    5264, 
    4636, 
    4723, 
    2552, 
    4708, 
    4438, 
    5887, 
    2591, 
    4438, 
    5693, 
    2591, 
    3600, 
    4438, 
    3938, 
    5771, 
    1249, 
    4428, 
    716, 
    1955, 
    1249, 
    5771, 
    1955, 
    1618, 
    787, 
    6193, 
    941, 
    1726, 
    1386, 
    6456, 
    2766, 
    5671, 
    1609, 
    5304, 
    774, 
    2449, 
    2766, 
    3129, 
    5692, 
    444, 
    443, 
    3661, 
    5692, 
    443, 
    3661, 
    1587, 
    5692, 
    6637, 
    413, 
    412, 
    411, 
    6637, 
    412, 
    411, 
    1258, 
    6637, 
    409, 
    755, 
    410, 
    6635, 
    391, 
    390, 
    641, 
    6635, 
    390, 
    6636, 
    392, 
    6635, 
    641, 
    6636, 
    6635, 
    641, 
    389, 
    6686, 
    6635, 
    392, 
    391, 
    641, 
    6686, 
    6636, 
    6686, 
    392, 
    6636, 
    2192, 
    6686, 
    389, 
    2192, 
    4670, 
    6686, 
    407, 
    4084, 
    408, 
    832, 
    1902, 
    405, 
    6654, 
    395, 
    394, 
    393, 
    2162, 
    5434, 
    6568, 
    400, 
    2300, 
    401, 
    6568, 
    402, 
    401, 
    400, 
    6568, 
    2091, 
    397, 
    2300, 
    398, 
    2091, 
    399, 
    398, 
    397, 
    2091, 
    399, 
    2091, 
    400, 
    400, 
    2091, 
    2300, 
    2300, 
    403, 
    402, 
    2300, 
    402, 
    6568, 
    1351, 
    2300, 
    397, 
    404, 
    403, 
    2300, 
    1351, 
    397, 
    396, 
    404, 
    1351, 
    405, 
    404, 
    2300, 
    1351, 
    5434, 
    2162, 
    1351, 
    6654, 
    5434, 
    396, 
    395, 
    6654, 
    396, 
    394, 
    5434, 
    6654, 
    394, 
    393, 
    5434, 
    5434, 
    1351, 
    396, 
    1090, 
    2162, 
    393, 
    1090, 
    832, 
    2162, 
    1351, 
    2162, 
    405, 
    1902, 
    642, 
    406, 
    405, 
    1902, 
    406, 
    2019, 
    407, 
    642, 
    832, 
    2019, 
    1902, 
    832, 
    4185, 
    2361, 
    2162, 
    832, 
    405, 
    392, 
    6686, 
    4670, 
    389, 
    388, 
    1167, 
    4084, 
    984, 
    409, 
    2019, 
    4084, 
    407, 
    2361, 
    5362, 
    4084, 
    832, 
    2361, 
    2019, 
    5362, 
    726, 
    984, 
    1878, 
    5362, 
    2361, 
    1878, 
    2302, 
    5362, 
    2019, 
    642, 
    1902, 
    1141, 
    1878, 
    4185, 
    1167, 
    388, 
    6619, 
    1076, 
    1994, 
    386, 
    2192, 
    389, 
    1167, 
    1141, 
    2192, 
    1167, 
    1141, 
    4185, 
    4670, 
    6619, 
    386, 
    1994, 
    387, 
    6619, 
    388, 
    387, 
    386, 
    6619, 
    1994, 
    1167, 
    6619, 
    1312, 
    1994, 
    1076, 
    1312, 
    1167, 
    1994, 
    1121, 
    385, 
    384, 
    3199, 
    726, 
    1284, 
    1301, 
    3199, 
    938, 
    984, 
    726, 
    3199, 
    408, 
    4084, 
    409, 
    4084, 
    2019, 
    2361, 
    4461, 
    385, 
    1121, 
    1284, 
    2302, 
    1442, 
    938, 
    1284, 
    771, 
    2302, 
    1878, 
    1141, 
    1442, 
    2302, 
    1312, 
    726, 
    5362, 
    2302, 
    386, 
    385, 
    1076, 
    984, 
    755, 
    409, 
    5761, 
    1740, 
    954, 
    2126, 
    4361, 
    1030, 
    1053, 
    1740, 
    4361, 
    2874, 
    3568, 
    1390, 
    4849, 
    1379, 
    1458, 
    2390, 
    4849, 
    1458, 
    1360, 
    2335, 
    4849, 
    4849, 
    2335, 
    1379, 
    4989, 
    1133, 
    1871, 
    4882, 
    4906, 
    2126, 
    5283, 
    4340, 
    1606, 
    4882, 
    5034, 
    4906, 
    4882, 
    3164, 
    5034, 
    5283, 
    5034, 
    4340, 
    1133, 
    5283, 
    1606, 
    1133, 
    4906, 
    5283, 
    1030, 
    4882, 
    2126, 
    1030, 
    3483, 
    4882, 
    1442, 
    1606, 
    771, 
    1442, 
    1076, 
    4461, 
    6062, 
    2377, 
    674, 
    1533, 
    6062, 
    674, 
    4989, 
    1871, 
    6062, 
    1121, 
    1871, 
    1133, 
    1121, 
    383, 
    1871, 
    2042, 
    878, 
    1663, 
    3568, 
    3842, 
    1390, 
    3842, 
    3109, 
    2042, 
    1390, 
    3842, 
    2042, 
    954, 
    1740, 
    3842, 
    3260, 
    5761, 
    954, 
    3109, 
    878, 
    2042, 
    1053, 
    3109, 
    1740, 
    1053, 
    1285, 
    3697, 
    2126, 
    1053, 
    4361, 
    1549, 
    701, 
    4573, 
    4195, 
    1549, 
    1285, 
    1053, 
    4195, 
    1285, 
    1533, 
    674, 
    4195, 
    4195, 
    4322, 
    1549, 
    1207, 
    1184, 
    2217, 
    2189, 
    1619, 
    1207, 
    1556, 
    2189, 
    1137, 
    1556, 
    714, 
    2189, 
    1619, 
    789, 
    1925, 
    2217, 
    2231, 
    1207, 
    714, 
    1780, 
    1619, 
    782, 
    6199, 
    1301, 
    5383, 
    3769, 
    2335, 
    3137, 
    5383, 
    2777, 
    5289, 
    3769, 
    5383, 
    6343, 
    5289, 
    5383, 
    6199, 
    6343, 
    3461, 
    6199, 
    5289, 
    6343, 
    3164, 
    3769, 
    5289, 
    2777, 
    842, 
    5634, 
    5612, 
    3137, 
    5634, 
    6199, 
    3461, 
    3414, 
    2810, 
    3164, 
    5289, 
    2023, 
    2777, 
    1360, 
    5612, 
    6523, 
    6281, 
    5634, 
    2711, 
    5612, 
    2777, 
    5634, 
    3137, 
    3087, 
    2711, 
    5634, 
    1657, 
    3087, 
    842, 
    4238, 
    2217, 
    3667, 
    3414, 
    6281, 
    1258, 
    6523, 
    3133, 
    6281, 
    2711, 
    6523, 
    5612, 
    3746, 
    3133, 
    6523, 
    1208, 
    742, 
    3133, 
    413, 
    6637, 
    1258, 
    1301, 
    755, 
    3199, 
    384, 
    383, 
    1121, 
    4195, 
    674, 
    4322, 
    2126, 
    1533, 
    4195, 
    3164, 
    4340, 
    5034, 
    4906, 
    4989, 
    2126, 
    6062, 
    1871, 
    2377, 
    2126, 
    4989, 
    1533, 
    4906, 
    1133, 
    4989, 
    4461, 
    1121, 
    1133, 
    1606, 
    4461, 
    1133, 
    1076, 
    385, 
    4461, 
    6705, 
    381, 
    2377, 
    383, 
    6705, 
    2377, 
    383, 
    382, 
    6705, 
    382, 
    381, 
    6705, 
    1650, 
    826, 
    673, 
    2211, 
    1650, 
    1933, 
    1170, 
    2211, 
    1219, 
    3628, 
    2611, 
    2668, 
    4733, 
    3628, 
    3896, 
    2211, 
    4733, 
    2787, 
    1170, 
    3628, 
    4733, 
    1170, 
    1899, 
    3628, 
    5026, 
    1502, 
    1063, 
    5026, 
    4874, 
    3467, 
    1820, 
    5026, 
    1063, 
    6104, 
    1191, 
    3812, 
    1820, 
    5889, 
    5026, 
    1820, 
    1191, 
    5889, 
    3145, 
    3896, 
    3467, 
    6104, 
    5889, 
    1191, 
    3145, 
    4733, 
    3896, 
    2211, 
    2787, 
    1650, 
    2211, 
    1170, 
    4733, 
    2390, 
    866, 
    4849, 
    1820, 
    2390, 
    1458, 
    1875, 
    866, 
    2390, 
    4399, 
    1875, 
    1063, 
    1502, 
    4399, 
    1063, 
    1502, 
    1556, 
    4399, 
    1137, 
    1677, 
    1875, 
    1925, 
    1184, 
    1207, 
    1619, 
    1925, 
    1207, 
    789, 
    1998, 
    4384, 
    1677, 
    866, 
    1875, 
    2231, 
    1677, 
    1137, 
    842, 
    866, 
    1677, 
    4167, 
    701, 
    1590, 
    1036, 
    1802, 
    671, 
    1684, 
    849, 
    878, 
    2339, 
    1365, 
    1217, 
    1931, 
    2339, 
    1217, 
    4413, 
    1519, 
    1359, 
    1802, 
    4413, 
    2339, 
    1802, 
    2811, 
    4413, 
    3434, 
    5825, 
    3105, 
    1365, 
    3422, 
    2029, 
    1018, 
    1791, 
    3422, 
    3109, 
    3842, 
    1740, 
    849, 
    1663, 
    878, 
    3568, 
    1458, 
    1379, 
    1191, 
    2874, 
    1390, 
    1191, 
    1820, 
    2874, 
    4703, 
    2787, 
    3145, 
    4849, 
    866, 
    2023, 
    2390, 
    1063, 
    1875, 
    3568, 
    2874, 
    1458, 
    954, 
    3568, 
    1379, 
    954, 
    3842, 
    3568, 
    1820, 
    1063, 
    2390, 
    2874, 
    1820, 
    1458, 
    6104, 
    3812, 
    6094, 
    4703, 
    6104, 
    6094, 
    4874, 
    5889, 
    6104, 
    4874, 
    5026, 
    5889, 
    3145, 
    4874, 
    4703, 
    3467, 
    1502, 
    5026, 
    1933, 
    1219, 
    2211, 
    673, 
    1933, 
    1650, 
    6206, 
    1532, 
    1344, 
    6206, 
    3857, 
    1532, 
    6011, 
    6206, 
    1029, 
    6011, 
    3857, 
    6206, 
    3585, 
    2707, 
    3857, 
    1686, 
    880, 
    2409, 
    4399, 
    1137, 
    1875, 
    4340, 
    782, 
    771, 
    1606, 
    4340, 
    771, 
    3164, 
    3483, 
    3769, 
    4361, 
    5761, 
    1030, 
    5383, 
    1360, 
    2777, 
    3260, 
    2335, 
    1796, 
    6343, 
    5383, 
    3137, 
    3260, 
    1379, 
    2335, 
    5761, 
    3260, 
    1796, 
    1030, 
    5761, 
    1796, 
    4361, 
    1740, 
    5761, 
    954, 
    1379, 
    3260, 
    2023, 
    842, 
    2777, 
    4849, 
    2023, 
    1360, 
    842, 
    3087, 
    5634, 
    3697, 
    3109, 
    1053, 
    4989, 
    6062, 
    1533, 
    383, 
    2377, 
    1871, 
    381, 
    1934, 
    2377, 
    5356, 
    380, 
    3816, 
    2377, 
    1934, 
    674, 
    381, 
    380, 
    1934, 
    3816, 
    378, 
    1239, 
    1590, 
    3816, 
    1239, 
    380, 
    379, 
    3816, 
    1067, 
    439, 
    438, 
    1067, 
    792, 
    646, 
    437, 
    1067, 
    438, 
    3550, 
    1054, 
    2141, 
    792, 
    3550, 
    2141, 
    1240, 
    2481, 
    3550, 
    437, 
    1240, 
    1067, 
    2254, 
    645, 
    1702, 
    439, 
    1067, 
    646, 
    6634, 
    441, 
    440, 
    792, 
    440, 
    646, 
    6634, 
    440, 
    702, 
    442, 
    6634, 
    702, 
    442, 
    441, 
    6634, 
    792, 
    702, 
    440, 
    2481, 
    2254, 
    4432, 
    1054, 
    2481, 
    1813, 
    1054, 
    3550, 
    2481, 
    6485, 
    644, 
    436, 
    1020, 
    1769, 
    988, 
    5927, 
    2506, 
    1497, 
    999, 
    5927, 
    1020, 
    2782, 
    2506, 
    5927, 
    1777, 
    2897, 
    999, 
    2345, 
    1380, 
    2782, 
    1315, 
    1998, 
    1331, 
    2305, 
    1521, 
    1315, 
    1998, 
    1248, 
    1331, 
    1521, 
    4384, 
    1315, 
    789, 
    1248, 
    1998, 
    645, 
    644, 
    906, 
    5844, 
    6485, 
    5202, 
    2878, 
    434, 
    433, 
    4684, 
    5006, 
    1840, 
    6006, 
    434, 
    2362, 
    1240, 
    792, 
    1067, 
    906, 
    3353, 
    1702, 
    6488, 
    1153, 
    1419, 
    3555, 
    5473, 
    3244, 
    2903, 
    1101, 
    1850, 
    2834, 
    6151, 
    5065, 
    3244, 
    5473, 
    6253, 
    2488, 
    1850, 
    1101, 
    1172, 
    5409, 
    1101, 
    1346, 
    2637, 
    2488, 
    1346, 
    1777, 
    2637, 
    1054, 
    1346, 
    1327, 
    2637, 
    1153, 
    1850, 
    2488, 
    2637, 
    1850, 
    1777, 
    999, 
    6316, 
    2897, 
    2782, 
    999, 
    1346, 
    2897, 
    1777, 
    1813, 
    2345, 
    2897, 
    3020, 
    1380, 
    2345, 
    1813, 
    6054, 
    2345, 
    6485, 
    435, 
    5202, 
    906, 
    6485, 
    5844, 
    436, 
    435, 
    6485, 
    6006, 
    2362, 
    5006, 
    5622, 
    6006, 
    5006, 
    5202, 
    435, 
    6006, 
    3020, 
    5844, 
    5074, 
    435, 
    434, 
    6006, 
    5622, 
    5074, 
    6006, 
    5927, 
    1497, 
    1020, 
    2918, 
    2506, 
    2782, 
    2037, 
    2918, 
    1380, 
    2037, 
    5418, 
    2918, 
    5418, 
    867, 
    3943, 
    3020, 
    5074, 
    1380, 
    5899, 
    1907, 
    1521, 
    2918, 
    5418, 
    2506, 
    3943, 
    1678, 
    3373, 
    6316, 
    1419, 
    1153, 
    1020, 
    3752, 
    999, 
    988, 
    1419, 
    3752, 
    4384, 
    1907, 
    1925, 
    789, 
    4384, 
    1925, 
    1998, 
    1315, 
    4384, 
    5232, 
    1769, 
    1020, 
    1521, 
    5232, 
    1497, 
    2305, 
    1769, 
    5232, 
    1711, 
    2305, 
    1315, 
    1711, 
    808, 
    2305, 
    5899, 
    2506, 
    5418, 
    1907, 
    5899, 
    2567, 
    1497, 
    2506, 
    5899, 
    999, 
    2782, 
    5927, 
    1907, 
    1184, 
    1925, 
    1497, 
    5899, 
    1521, 
    3943, 
    867, 
    1678, 
    2656, 
    6027, 
    3040, 
    5418, 
    2037, 
    867, 
    6144, 
    5418, 
    3943, 
    2567, 
    5899, 
    5418, 
    5908, 
    6488, 
    3351, 
    2878, 
    433, 
    432, 
    1840, 
    2878, 
    432, 
    2362, 
    434, 
    2878, 
    2232, 
    3373, 
    1678, 
    2656, 
    3667, 
    1184, 
    1907, 
    6027, 
    1184, 
    3746, 
    1208, 
    3133, 
    4585, 
    3746, 
    2711, 
    3373, 
    2232, 
    3746, 
    1657, 
    2231, 
    2217, 
    2217, 
    4238, 
    1657, 
    1184, 
    3667, 
    2217, 
    2656, 
    3040, 
    3667, 
    842, 
    1677, 
    1657, 
    1204, 
    1415, 
    424, 
    1204, 
    423, 
    422, 
    2427, 
    1415, 
    1204, 
    428, 
    2427, 
    813, 
    427, 
    426, 
    2427, 
    424, 
    423, 
    1204, 
    1415, 
    425, 
    424, 
    1638, 
    2427, 
    1204, 
    426, 
    425, 
    1415, 
    1638, 
    422, 
    2067, 
    2427, 
    1638, 
    813, 
    1204, 
    422, 
    1638, 
    426, 
    1415, 
    2427, 
    813, 
    429, 
    428, 
    427, 
    2427, 
    428, 
    2067, 
    421, 
    697, 
    1638, 
    2067, 
    1423, 
    422, 
    421, 
    2067, 
    1947, 
    2067, 
    697, 
    1947, 
    697, 
    5342, 
    430, 
    1947, 
    1376, 
    1423, 
    2067, 
    1947, 
    813, 
    1423, 
    429, 
    813, 
    1638, 
    1423, 
    1423, 
    430, 
    429, 
    420, 
    697, 
    421, 
    4779, 
    419, 
    418, 
    1427, 
    5342, 
    6347, 
    420, 
    419, 
    4779, 
    418, 
    1812, 
    4779, 
    417, 
    416, 
    6696, 
    823, 
    2373, 
    4828, 
    1427, 
    823, 
    1647, 
    1947, 
    5342, 
    1376, 
    4828, 
    416, 
    415, 
    823, 
    4828, 
    1342, 
    1812, 
    416, 
    4828, 
    6347, 
    4779, 
    1812, 
    2373, 
    6347, 
    1812, 
    5342, 
    4779, 
    6347, 
    1376, 
    5342, 
    1427, 
    697, 
    4779, 
    5342, 
    6696, 
    416, 
    1812, 
    418, 
    6696, 
    1812, 
    418, 
    417, 
    6696, 
    4828, 
    415, 
    1342, 
    924, 
    1376, 
    1427, 
    2960, 
    1576, 
    5119, 
    643, 
    2208, 
    976, 
    1647, 
    823, 
    1476, 
    2208, 
    1647, 
    1015, 
    924, 
    1427, 
    1647, 
    430, 
    924, 
    431, 
    4779, 
    697, 
    420, 
    430, 
    1376, 
    924, 
    430, 
    1423, 
    1947, 
    924, 
    2208, 
    431, 
    2373, 
    823, 
    1427, 
    6347, 
    2373, 
    1427, 
    1812, 
    4828, 
    2373, 
    2960, 
    1342, 
    415, 
    4317, 
    1208, 
    2232, 
    5119, 
    1576, 
    1476, 
    823, 
    5119, 
    1476, 
    1342, 
    2960, 
    5119, 
    742, 
    1208, 
    1576, 
    2208, 
    643, 
    431, 
    1647, 
    2208, 
    924, 
    1015, 
    976, 
    2208, 
    2960, 
    413, 
    742, 
    2960, 
    742, 
    1576, 
    414, 
    2960, 
    415, 
    414, 
    413, 
    2960, 
    6281, 
    3133, 
    413, 
    1258, 
    6281, 
    413, 
    3414, 
    5612, 
    6281, 
    1301, 
    3414, 
    1258, 
    6523, 
    2711, 
    3746, 
    3461, 
    5612, 
    3414, 
    3461, 
    3137, 
    5612, 
    4684, 
    1678, 
    867, 
    1476, 
    4317, 
    1091, 
    2232, 
    1678, 
    4064, 
    1091, 
    4317, 
    4064, 
    4585, 
    2711, 
    4238, 
    3040, 
    4585, 
    3667, 
    3040, 
    3373, 
    4585, 
    6027, 
    6144, 
    3040, 
    1184, 
    6027, 
    2656, 
    6144, 
    3943, 
    3040, 
    2567, 
    6144, 
    6027, 
    2567, 
    5418, 
    6144, 
    3373, 
    3746, 
    4585, 
    3943, 
    3373, 
    3040, 
    2232, 
    1208, 
    3746, 
    413, 
    3133, 
    742, 
    5074, 
    5622, 
    2037, 
    4064, 
    4684, 
    1840, 
    4064, 
    1678, 
    4684, 
    4238, 
    3087, 
    1657, 
    4585, 
    4238, 
    3667, 
    2711, 
    3087, 
    4238, 
    6027, 
    1907, 
    2567, 
    2231, 
    2189, 
    1207, 
    1677, 
    2231, 
    1657, 
    1137, 
    2189, 
    2231, 
    1907, 
    4384, 
    1521, 
    4777, 
    976, 
    1015, 
    6199, 
    782, 
    2810, 
    5289, 
    6199, 
    2810, 
    3414, 
    1301, 
    6199, 
    755, 
    1301, 
    1258, 
    938, 
    782, 
    1301, 
    984, 
    3199, 
    755, 
    3199, 
    1284, 
    938, 
    2722, 
    1359, 
    1018, 
    841, 
    1519, 
    2811, 
    5822, 
    4616, 
    2495, 
    5822, 
    4786, 
    4616, 
    3343, 
    5822, 
    3007, 
    6139, 
    1519, 
    841, 
    3343, 
    6139, 
    5822, 
    3343, 
    1359, 
    6139, 
    841, 
    1656, 
    4786, 
    4322, 
    701, 
    1549, 
    1934, 
    4322, 
    674, 
    1934, 
    5356, 
    4322, 
    2909, 
    2495, 
    4416, 
    1148, 
    2909, 
    890, 
    1148, 
    1885, 
    4377, 
    1663, 
    5067, 
    1390, 
    6206, 
    1344, 
    1029, 
    3147, 
    5960, 
    2789, 
    673, 
    826, 
    1532, 
    5067, 
    3535, 
    3812, 
    3697, 
    878, 
    3109, 
    1285, 
    4775, 
    3697, 
    2029, 
    849, 
    1684, 
    2236, 
    2029, 
    1684, 
    1365, 
    2722, 
    3422, 
    3816, 
    379, 
    378, 
    2727, 
    4080, 
    377, 
    4167, 
    5865, 
    1931, 
    1217, 
    4573, 
    1931, 
    1590, 
    1239, 
    5865, 
    4322, 
    5356, 
    701, 
    5865, 
    4080, 
    671, 
    1590, 
    5865, 
    4167, 
    1239, 
    4080, 
    5865, 
    5356, 
    3816, 
    1590, 
    701, 
    5356, 
    1590, 
    1934, 
    380, 
    5356, 
    378, 
    377, 
    1239, 
    755, 
    1258, 
    411, 
    410, 
    755, 
    411, 
    4195, 
    1053, 
    2126, 
    4775, 
    2236, 
    3697, 
    4573, 
    4775, 
    1549, 
    4573, 
    1217, 
    4775, 
    2236, 
    1365, 
    2029, 
    3697, 
    2236, 
    1684, 
    878, 
    3697, 
    1684, 
    1285, 
    1549, 
    4775, 
    1217, 
    1365, 
    2236, 
    3535, 
    5723, 
    2017, 
    3434, 
    3105, 
    5067, 
    3422, 
    3434, 
    849, 
    5825, 
    1791, 
    1029, 
    3422, 
    5825, 
    3434, 
    3422, 
    1791, 
    5825, 
    5825, 
    1029, 
    3105, 
    3769, 
    3483, 
    1796, 
    1360, 
    5383, 
    2335, 
    3137, 
    3461, 
    6343, 
    4340, 
    3164, 
    2810, 
    782, 
    4340, 
    2810, 
    5034, 
    5283, 
    4906, 
    3769, 
    1796, 
    2335, 
    4882, 
    3483, 
    3164, 
    1030, 
    1796, 
    3483, 
    2017, 
    5723, 
    1344, 
    826, 
    3535, 
    2017, 
    5067, 
    1663, 
    3434, 
    5723, 
    5067, 
    3105, 
    1344, 
    5723, 
    3105, 
    3535, 
    5067, 
    5723, 
    3812, 
    1390, 
    5067, 
    826, 
    1650, 
    6094, 
    1191, 
    1390, 
    3812, 
    2042, 
    1663, 
    1390, 
    849, 
    3434, 
    1663, 
    866, 
    842, 
    2023, 
    938, 
    771, 
    782, 
    4670, 
    1090, 
    393, 
    392, 
    4670, 
    393, 
    2192, 
    1141, 
    4670, 
    1312, 
    1141, 
    1167, 
    1442, 
    1312, 
    1076, 
    4461, 
    1606, 
    1442, 
    771, 
    1284, 
    1442, 
    1284, 
    726, 
    2302, 
    4185, 
    832, 
    1090, 
    4670, 
    4185, 
    1090, 
    1878, 
    2361, 
    4185, 
    1312, 
    2302, 
    1141, 
    5362, 
    984, 
    4084, 
    375, 
    374, 
    2124, 
    2131, 
    2124, 
    1205, 
    2189, 
    714, 
    1619, 
    4399, 
    1556, 
    1137, 
    5685, 
    3467, 
    3896, 
    2668, 
    5685, 
    3896, 
    3050, 
    1556, 
    5685, 
    6094, 
    3812, 
    3535, 
    826, 
    6094, 
    3535, 
    4703, 
    4874, 
    6104, 
    2787, 
    4703, 
    1650, 
    3145, 
    3467, 
    4874, 
    3628, 
    1899, 
    2611, 
    3668, 
    1618, 
    2188, 
    1135, 
    3668, 
    2188, 
    5294, 
    3828, 
    3555, 
    4046, 
    4753, 
    3110, 
    4094, 
    3828, 
    4753, 
    4312, 
    4094, 
    4046, 
    787, 
    4312, 
    4046, 
    1618, 
    3668, 
    4312, 
    6186, 
    3828, 
    4094, 
    5662, 
    6186, 
    4094, 
    3367, 
    3035, 
    6186, 
    1135, 
    3530, 
    3668, 
    6186, 
    5473, 
    3828, 
    5674, 
    3218, 
    2867, 
    3668, 
    4673, 
    3367, 
    3530, 
    3218, 
    4673, 
    3668, 
    3530, 
    4673, 
    1135, 
    1874, 
    3530, 
    6488, 
    5908, 
    2834, 
    1635, 
    6488, 
    1419, 
    1635, 
    3351, 
    6488, 
    6151, 
    3244, 
    5065, 
    5294, 
    6151, 
    3184, 
    3555, 
    3244, 
    6151, 
    3110, 
    4753, 
    5294, 
    6253, 
    2649, 
    4070, 
    3828, 
    5473, 
    3555, 
    3035, 
    2649, 
    5473, 
    3244, 
    2903, 
    5065, 
    3440, 
    5294, 
    3184, 
    6253, 
    4070, 
    6148, 
    2903, 
    6253, 
    6148, 
    5473, 
    2649, 
    6253, 
    6448, 
    6164, 
    5713, 
    5803, 
    6448, 
    5713, 
    5652, 
    2449, 
    6448, 
    5065, 
    1850, 
    1153, 
    3184, 
    6151, 
    2834, 
    2903, 
    1850, 
    5065, 
    6193, 
    4428, 
    1618, 
    3929, 
    6193, 
    787, 
    3929, 
    716, 
    6193, 
    2389, 
    4720, 
    1874, 
    4720, 
    3218, 
    3530, 
    1874, 
    4720, 
    3530, 
    5996, 
    6385, 
    3766, 
    5671, 
    5996, 
    3766, 
    5042, 
    4895, 
    6385, 
    2389, 
    4825, 
    4720, 
    2389, 
    1456, 
    4825, 
    3218, 
    5674, 
    4673, 
    5652, 
    6449, 
    2449, 
    5674, 
    3035, 
    4673, 
    2449, 
    6449, 
    2867, 
    6541, 
    5803, 
    4070, 
    2867, 
    6449, 
    5674, 
    5652, 
    5803, 
    6449, 
    4428, 
    2188, 
    1618, 
    3938, 
    1135, 
    2188, 
    5771, 
    3938, 
    2188, 
    4428, 
    5771, 
    2188, 
    4428, 
    1955, 
    5771, 
    1249, 
    2262, 
    3938, 
    923, 
    5569, 
    1222, 
    4343, 
    4622, 
    1557, 
    6046, 
    5788, 
    4131, 
    3868, 
    6046, 
    4131, 
    5828, 
    5682, 
    6046, 
    2146, 
    4343, 
    1557, 
    4035, 
    4131, 
    4343, 
    5828, 
    3598, 
    5611, 
    5505, 
    5611, 
    3294, 
    2955, 
    5505, 
    3294, 
    3988, 
    4215, 
    5492, 
    2146, 
    4035, 
    4343, 
    5172, 
    1065, 
    1822, 
    5036, 
    5172, 
    3443, 
    5036, 
    4259, 
    5172, 
    4131, 
    4035, 
    4259, 
    2146, 
    1065, 
    4035, 
    5583, 
    5618, 
    2550, 
    5828, 
    3868, 
    3598, 
    5934, 
    5828, 
    5611, 
    5721, 
    5934, 
    5611, 
    5543, 
    5800, 
    5934, 
    5682, 
    6303, 
    6046, 
    5934, 
    5800, 
    5682, 
    6303, 
    4215, 
    4429, 
    6046, 
    6303, 
    5788, 
    5492, 
    4215, 
    6303, 
    5611, 
    3598, 
    3294, 
    5721, 
    5611, 
    5505, 
    5800, 
    5644, 
    5682, 
    5828, 
    5934, 
    5682, 
    5543, 
    6200, 
    5800, 
    3809, 
    3498, 
    3532, 
    4833, 
    2923, 
    2512, 
    3369, 
    6344, 
    3037, 
    4477, 
    3265, 
    4657, 
    4268, 
    6239, 
    5564, 
    5564, 
    3573, 
    3265, 
    4477, 
    5564, 
    3265, 
    4477, 
    4268, 
    5564, 
    2869, 
    4268, 
    2451, 
    4042, 
    6135, 
    6239, 
    6272, 
    4371, 
    4522, 
    3179, 
    6272, 
    5754, 
    3179, 
    2828, 
    6272, 
    6480, 
    6262, 
    5620, 
    5657, 
    6480, 
    5835, 
    6349, 
    6262, 
    6480, 
    6353, 
    6452, 
    6519, 
    6293, 
    6262, 
    6349, 
    5864, 
    6203, 
    6464, 
    6203, 
    4326, 
    6329, 
    4371, 
    6115, 
    6086, 
    5689, 
    5499, 
    5810, 
    5835, 
    5689, 
    5657, 
    6349, 
    6480, 
    5657, 
    5620, 
    5511, 
    5835, 
    6160, 
    5547, 
    5751, 
    5689, 
    6042, 
    5499, 
    5696, 
    5547, 
    6042, 
    5511, 
    5696, 
    5689, 
    5511, 
    6001, 
    6137, 
    6549, 
    6564, 
    6416, 
    5750, 
    6549, 
    6416, 
    6434, 
    3885, 
    6564, 
    5864, 
    3845, 
    4112, 
    5864, 
    5470, 
    3845, 
    4326, 
    6203, 
    4112, 
    5724, 
    5470, 
    5864, 
    6262, 
    6086, 
    5620, 
    6464, 
    5724, 
    5864, 
    6349, 
    6562, 
    6293, 
    6426, 
    5724, 
    6464, 
    6293, 
    6329, 
    6262, 
    4112, 
    6203, 
    5864, 
    6329, 
    6086, 
    6262, 
    6203, 
    6329, 
    6293, 
    4326, 
    4522, 
    6329, 
    5724, 
    6208, 
    5779, 
    6375, 
    5945, 
    5784, 
    5689, 
    5810, 
    5657, 
    6366, 
    6040, 
    5914, 
    5780, 
    6417, 
    5914, 
    6543, 
    6364, 
    6481, 
    6560, 
    6543, 
    6376, 
    6490, 
    6560, 
    6376, 
    6565, 
    6559, 
    6543, 
    6540, 
    6565, 
    6560, 
    6540, 
    6539, 
    6565, 
    6565, 
    6539, 
    6559, 
    6543, 
    6560, 
    6565, 
    6490, 
    6366, 
    6560, 
    6366, 
    6461, 
    6540, 
    6365, 
    6482, 
    6539, 
    5499, 
    5945, 
    5810, 
    6158, 
    6376, 
    6377, 
    5705, 
    5829, 
    5483, 
    6096, 
    5683, 
    5518, 
    6459, 
    6028, 
    5765, 
    5748, 
    5559, 
    5651, 
    6275, 
    6178, 
    5748, 
    6338, 
    6275, 
    5581, 
    5904, 
    6338, 
    5581, 
    5617, 
    6089, 
    6338, 
    6483, 
    5841, 
    6462, 
    5979, 
    6483, 
    6275, 
    5979, 
    5841, 
    6483, 
    6474, 
    5804, 
    4351, 
    6064, 
    5938, 
    6465, 
    6178, 
    6064, 
    6467, 
    5581, 
    6275, 
    5748, 
    6275, 
    6483, 
    6178, 
    6512, 
    5695, 
    5509, 
    5938, 
    6512, 
    6416, 
    6462, 
    5695, 
    6512, 
    6178, 
    6462, 
    6064, 
    6178, 
    6483, 
    6462, 
    6064, 
    6462, 
    6512, 
    5735, 
    4964, 
    4723, 
    6467, 
    6064, 
    6465, 
    5748, 
    6467, 
    5559, 
    5748, 
    6178, 
    6467, 
    5938, 
    6064, 
    6512, 
    6416, 
    6564, 
    5804, 
    6474, 
    4351, 
    2591, 
    6465, 
    6474, 
    4964, 
    6465, 
    5938, 
    6474, 
    6416, 
    5804, 
    5938, 
    5750, 
    6416, 
    5509, 
    6549, 
    5583, 
    6434, 
    4140, 
    4351, 
    5804, 
    4636, 
    6457, 
    4723, 
    5035, 
    3369, 
    4419, 
    4618, 
    5035, 
    4419, 
    4883, 
    2869, 
    5035, 
    4880, 
    4536, 
    1874, 
    2262, 
    4880, 
    3938, 
    2262, 
    1712, 
    4880, 
    2141, 
    1327, 
    828, 
    1240, 
    3550, 
    792, 
    1054, 
    1327, 
    2141, 
    828, 
    3661, 
    443, 
    1327, 
    5409, 
    828, 
    3367, 
    4673, 
    3035, 
    1346, 
    2488, 
    1327, 
    6316, 
    1153, 
    2637, 
    1777, 
    6316, 
    2637, 
    3752, 
    1419, 
    6316, 
    1769, 
    1635, 
    988, 
    3927, 
    4576, 
    4751, 
    4046, 
    4094, 
    4753, 
    1997, 
    4046, 
    2743, 
    787, 
    1618, 
    4312, 
    5699, 
    3351, 
    2728, 
    3719, 
    5699, 
    2728, 
    3719, 
    3655, 
    5699, 
    3927, 
    3655, 
    3719, 
    3100, 
    3927, 
    3428, 
    5772, 
    3440, 
    3184, 
    3927, 
    4751, 
    3655, 
    6061, 
    3440, 
    5772, 
    4576, 
    6061, 
    4751, 
    4576, 
    3110, 
    6061, 
    5908, 
    3184, 
    2834, 
    4751, 
    5772, 
    3655, 
    4751, 
    6061, 
    5772, 
    5294, 
    3555, 
    6151, 
    3110, 
    5294, 
    3440, 
    4753, 
    3828, 
    5294, 
    2743, 
    4046, 
    3110, 
    6186, 
    3035, 
    5473, 
    5772, 
    5908, 
    3655, 
    988, 
    1635, 
    1419, 
    4576, 
    4169, 
    4382, 
    1153, 
    2834, 
    5065, 
    3668, 
    5662, 
    4312, 
    5692, 
    1587, 
    753, 
    5409, 
    3661, 
    828, 
    1172, 
    1587, 
    3661, 
    442, 
    702, 
    443, 
    6326, 
    3915, 
    3645, 
    2757, 
    6210, 
    2534, 
    6091, 
    4376, 
    5522, 
    4821, 
    6091, 
    5522, 
    4821, 
    4645, 
    6091, 
    4742, 
    4254, 
    4271, 
    5852, 
    4464, 
    4742, 
    4163, 
    5522, 
    4376, 
    5323, 
    2558, 
    5371, 
    4645, 
    5323, 
    5226, 
    4821, 
    6210, 
    5323, 
    6321, 
    2679, 
    2478, 
    5312, 
    6321, 
    4626, 
    5312, 
    2679, 
    6321, 
    4436, 
    5312, 
    4626, 
    5210, 
    5229, 
    5312, 
    4957, 
    5174, 
    5038, 
    5097, 
    5226, 
    5271, 
    4163, 
    5523, 
    2937, 
    5174, 
    4957, 
    5097, 
    4222, 
    5084, 
    5210, 
    4890, 
    4803, 
    5038, 
    1219, 
    2779, 
    2238, 
    1219, 
    1933, 
    4028, 
    2238, 
    1170, 
    1219, 
    4047, 
    673, 
    3083, 
    1686, 
    1899, 
    2238, 
    5376, 
    4254, 
    4464, 
    4645, 
    5376, 
    4464, 
    5097, 
    4957, 
    5452, 
    880, 
    5167, 
    2409, 
    5056, 
    1767, 
    4914, 
    1065, 
    5056, 
    1822, 
    2304, 
    1767, 
    5056, 
    2936, 
    2304, 
    5056, 
    2146, 
    2936, 
    1065, 
    1314, 
    2304, 
    2936, 
    4382, 
    4169, 
    2304, 
    2743, 
    4382, 
    1314, 
    2743, 
    3110, 
    4382, 
    2146, 
    4540, 
    2936, 
    5908, 
    5772, 
    3184, 
    1153, 
    6488, 
    2834, 
    3351, 
    3655, 
    5908, 
    808, 
    3351, 
    1635, 
    4169, 
    3100, 
    1767, 
    1314, 
    4382, 
    2304, 
    3927, 
    3100, 
    4169, 
    3719, 
    3428, 
    3927, 
    3351, 
    5699, 
    3655, 
    6198, 
    6166, 
    5410, 
    5647, 
    6198, 
    5410, 
    3719, 
    2728, 
    6198, 
    5410, 
    2491, 
    2723, 
    5647, 
    5410, 
    3716, 
    6198, 
    2728, 
    6166, 
    1997, 
    2743, 
    1314, 
    1997, 
    787, 
    4046, 
    5232, 
    1521, 
    2305, 
    1619, 
    1780, 
    789, 
    1769, 
    808, 
    1635, 
    1497, 
    5232, 
    1020, 
    2305, 
    808, 
    1769, 
    1331, 
    1711, 
    1315, 
    1331, 
    2491, 
    6166, 
    6433, 
    2723, 
    2491, 
    1780, 
    5575, 
    6433, 
    1780, 
    3641, 
    5575, 
    6166, 
    2728, 
    1711, 
    1331, 
    6166, 
    1711, 
    2491, 
    5410, 
    6166, 
    6155, 
    2723, 
    5575, 
    3715, 
    6155, 
    3335, 
    3715, 
    3423, 
    6155, 
    986, 
    5212, 
    2105, 
    6198, 
    3428, 
    3719, 
    5212, 
    5647, 
    3716, 
    5212, 
    3100, 
    5647, 
    6433, 
    5575, 
    2723, 
    1248, 
    6433, 
    1331, 
    1248, 
    1780, 
    6433, 
    3100, 
    986, 
    1767, 
    3420, 
    2105, 
    1485, 
    5167, 
    3420, 
    1485, 
    2044, 
    1391, 
    3420, 
    2906, 
    986, 
    2105, 
    3420, 
    2906, 
    2105, 
    1391, 
    2352, 
    2906, 
    2418, 
    2528, 
    1912, 
    4799, 
    6174, 
    4626, 
    4467, 
    3598, 
    3868, 
    4890, 
    4970, 
    880, 
    3114, 
    3994, 
    2747, 
    3730, 
    1391, 
    4944, 
    4436, 
    4211, 
    4222, 
    5662, 
    3367, 
    6186, 
    4312, 
    5662, 
    4094, 
    3668, 
    3367, 
    5662, 
    4540, 
    1997, 
    1314, 
    2936, 
    4540, 
    1314, 
    2146, 
    1557, 
    4540, 
    3929, 
    787, 
    1997, 
    4540, 
    3929, 
    1997, 
    1557, 
    716, 
    3929, 
    2728, 
    808, 
    1711, 
    3716, 
    3423, 
    5212, 
    3428, 
    6198, 
    5647, 
    2723, 
    6155, 
    3716, 
    6061, 
    3110, 
    3440, 
    4169, 
    4576, 
    3927, 
    4382, 
    3110, 
    4576, 
    5410, 
    2723, 
    3716, 
    1767, 
    2304, 
    4169, 
    2906, 
    2352, 
    4914, 
    2728, 
    3351, 
    808, 
    1780, 
    1248, 
    789, 
    4733, 
    3145, 
    2787, 
    2668, 
    3896, 
    3628, 
    2668, 
    3050, 
    5685, 
    5575, 
    3335, 
    6155, 
    3050, 
    3641, 
    1780, 
    3050, 
    2668, 
    3641, 
    5167, 
    1485, 
    2409, 
    2044, 
    5167, 
    880, 
    2044, 
    3420, 
    5167, 
    1686, 
    2238, 
    4803, 
    1391, 
    2906, 
    3420, 
    5212, 
    986, 
    3100, 
    3428, 
    5647, 
    3100, 
    3423, 
    2105, 
    5212, 
    2254, 
    1240, 
    437, 
    645, 
    2254, 
    437, 
    1702, 
    4432, 
    2254, 
    906, 
    1702, 
    645, 
    6054, 
    3353, 
    3020, 
    2345, 
    6054, 
    3020, 
    4432, 
    1702, 
    6054, 
    6485, 
    906, 
    644, 
    5074, 
    5844, 
    5202, 
    3353, 
    906, 
    5844, 
    976, 
    1840, 
    432, 
    976, 
    1091, 
    1840, 
    643, 
    976, 
    432, 
    5119, 
    823, 
    1342, 
    4317, 
    1476, 
    1576, 
    1208, 
    4317, 
    1576, 
    2232, 
    4064, 
    4317, 
    4777, 
    1015, 
    1476, 
    1091, 
    4777, 
    1476, 
    1091, 
    976, 
    4777, 
    1840, 
    1091, 
    4064, 
    5006, 
    2362, 
    1840, 
    867, 
    2037, 
    5622, 
    5844, 
    3020, 
    3353, 
    6006, 
    5074, 
    5202, 
    4684, 
    5622, 
    5006, 
    4684, 
    867, 
    5622, 
    2037, 
    1380, 
    5074, 
    2362, 
    2878, 
    1840, 
    1015, 
    1647, 
    1476, 
    3752, 
    1020, 
    988, 
    4080, 
    1530, 
    671, 
    376, 
    2727, 
    377, 
    376, 
    2124, 
    2727, 
    374, 
    373, 
    681, 
    372, 
    681, 
    373, 
    4851, 
    703, 
    834, 
    1653, 
    4931, 
    834, 
    2363, 
    1409, 
    4851, 
    3396, 
    4018, 
    1629, 
    800, 
    3691, 
    1629, 
    3065, 
    5494, 
    4018, 
    4055, 
    366, 
    365, 
    1409, 
    2880, 
    2058, 
    1241, 
    366, 
    2462, 
    4055, 
    908, 
    5308, 
    366, 
    4055, 
    2462, 
    365, 
    364, 
    4055, 
    2745, 
    5550, 
    1023, 
    2254, 
    2481, 
    1240, 
    4432, 
    1813, 
    2481, 
    3353, 
    6054, 
    1702, 
    6054, 
    1813, 
    4432, 
    2918, 
    2782, 
    1380, 
    2782, 
    2897, 
    2345, 
    2897, 
    1054, 
    1813, 
    3752, 
    6316, 
    999, 
    1346, 
    1054, 
    2897, 
    5409, 
    1327, 
    2488, 
    1101, 
    5409, 
    2488, 
    1172, 
    3661, 
    5409, 
    828, 
    702, 
    2141, 
    702, 
    792, 
    2141, 
    3050, 
    1780, 
    714, 
    3335, 
    2611, 
    2999, 
    3641, 
    2668, 
    3335, 
    1556, 
    3050, 
    714, 
    1556, 
    1502, 
    5685, 
    5685, 
    1502, 
    3467, 
    1899, 
    2409, 
    2611, 
    2238, 
    1899, 
    1170, 
    2409, 
    1485, 
    3715, 
    1686, 
    2409, 
    1899, 
    6433, 
    2491, 
    1331, 
    3641, 
    3335, 
    5575, 
    2611, 
    3335, 
    2668, 
    6155, 
    3423, 
    3716, 
    2999, 
    3715, 
    3335, 
    2999, 
    2409, 
    3715, 
    2409, 
    2999, 
    2611, 
    1485, 
    3423, 
    3715, 
    1485, 
    2105, 
    3423, 
    753, 
    445, 
    444, 
    702, 
    828, 
    443, 
    3766, 
    6385, 
    3480, 
    3218, 
    4895, 
    2867, 
    3218, 
    4720, 
    4895, 
    444, 
    5692, 
    753, 
    6148, 
    1101, 
    2903, 
    567, 
    566, 
    6622, 
    6622, 
    569, 
    568, 
    567, 
    6622, 
    568, 
    566, 
    6655, 
    6622, 
    6655, 
    569, 
    6622, 
    6624, 
    6655, 
    566, 
    6624, 
    569, 
    6655, 
    565, 
    6624, 
    566, 
    565, 
    6623, 
    6624, 
    6623, 
    565, 
    564, 
    569, 
    6623, 
    570, 
    569, 
    6624, 
    6623, 
    6656, 
    6623, 
    564, 
    2411, 
    6656, 
    564, 
    570, 
    6623, 
    6656, 
    2411, 
    570, 
    6656, 
    6682, 
    660, 
    6640, 
    563, 
    6682, 
    661, 
    563, 
    660, 
    6682, 
    660, 
    562, 
    6640, 
    6639, 
    562, 
    3577, 
    661, 
    6640, 
    564, 
    6640, 
    562, 
    6639, 
    564, 
    6640, 
    6639, 
    661, 
    6682, 
    6640, 
    6300, 
    562, 
    1038, 
    2411, 
    3577, 
    1489, 
    2411, 
    564, 
    3577, 
    560, 
    1349, 
    1473, 
    6666, 
    560, 
    559, 
    558, 
    6666, 
    559, 
    558, 
    1349, 
    6666, 
    6641, 
    658, 
    556, 
    555, 
    6641, 
    556, 
    555, 
    657, 
    6657, 
    555, 
    6657, 
    6641, 
    6704, 
    6626, 
    659, 
    658, 
    6704, 
    659, 
    6657, 
    657, 
    6704, 
    6641, 
    6657, 
    658, 
    657, 
    6626, 
    6704, 
    657, 
    554, 
    6626, 
    6626, 
    554, 
    1123, 
    557, 
    6626, 
    1123, 
    6704, 
    658, 
    6657, 
    1123, 
    554, 
    553, 
    2249, 
    553, 
    552, 
    557, 
    1123, 
    897, 
    557, 
    659, 
    6626, 
    2249, 
    897, 
    1123, 
    553, 
    2249, 
    1123, 
    552, 
    551, 
    2249, 
    897, 
    558, 
    557, 
    551, 
    964, 
    2249, 
    551, 
    550, 
    964, 
    2402, 
    831, 
    3852, 
    897, 
    1775, 
    1349, 
    964, 
    2314, 
    1775, 
    2249, 
    964, 
    897, 
    2314, 
    831, 
    1775, 
    550, 
    2314, 
    964, 
    550, 
    1325, 
    2314, 
    897, 
    964, 
    1775, 
    1325, 
    549, 
    548, 
    547, 
    5002, 
    548, 
    546, 
    4702, 
    547, 
    810, 
    4331, 
    1175, 
    1604, 
    2402, 
    3852, 
    2402, 
    1473, 
    1349, 
    5087, 
    1949, 
    707, 
    4526, 
    5087, 
    1604, 
    4526, 
    1949, 
    5087, 
    1986, 
    6020, 
    767, 
    1242, 
    1949, 
    4526, 
    2325, 
    1473, 
    1604, 
    5087, 
    2325, 
    1604, 
    707, 
    6300, 
    2325, 
    558, 
    897, 
    1349, 
    3254, 
    548, 
    5002, 
    2314, 
    1325, 
    831, 
    550, 
    549, 
    1325, 
    544, 
    6584, 
    545, 
    6584, 
    810, 
    4702, 
    6584, 
    656, 
    545, 
    810, 
    6584, 
    544, 
    4702, 
    656, 
    6584, 
    5427, 
    970, 
    4986, 
    5077, 
    1470, 
    1911, 
    1761, 
    5077, 
    4494, 
    1761, 
    2297, 
    5077, 
    1470, 
    861, 
    4598, 
    5002, 
    2200, 
    3254, 
    1175, 
    5002, 
    547, 
    1175, 
    2200, 
    5002, 
    4533, 
    1155, 
    2200, 
    1986, 
    4533, 
    851, 
    1986, 
    1155, 
    4533, 
    831, 
    1325, 
    3254, 
    4702, 
    546, 
    656, 
    1175, 
    4702, 
    810, 
    1175, 
    547, 
    4702, 
    4877, 
    1175, 
    4331, 
    4533, 
    2200, 
    4877, 
    3254, 
    1325, 
    548, 
    1155, 
    3254, 
    2200, 
    1155, 
    831, 
    3254, 
    5320, 
    2519, 
    1489, 
    4697, 
    5320, 
    2107, 
    4697, 
    4524, 
    5320, 
    6116, 
    4524, 
    4697, 
    4521, 
    6116, 
    4324, 
    4521, 
    5159, 
    6116, 
    1867, 
    2519, 
    4524, 
    571, 
    2411, 
    1445, 
    4484, 
    6300, 
    707, 
    6666, 
    1349, 
    560, 
    846, 
    1742, 
    1660, 
    6577, 
    539, 
    6578, 
    540, 
    6577, 
    541, 
    540, 
    539, 
    6577, 
    6578, 
    538, 
    537, 
    1675, 
    6579, 
    537, 
    539, 
    538, 
    6578, 
    6578, 
    6579, 
    6577, 
    6579, 
    541, 
    6577, 
    537, 
    6579, 
    6578, 
    1675, 
    541, 
    6579, 
    536, 
    1675, 
    537, 
    536, 
    1713, 
    1675, 
    655, 
    541, 
    1675, 
    1675, 
    920, 
    655, 
    2214, 
    836, 
    1761, 
    1179, 
    2214, 
    977, 
    1713, 
    836, 
    2214, 
    1675, 
    1713, 
    920, 
    535, 
    836, 
    1713, 
    1179, 
    920, 
    2214, 
    655, 
    920, 
    542, 
    536, 
    535, 
    1713, 
    535, 
    534, 
    836, 
    2214, 
    920, 
    1713, 
    2008, 
    1179, 
    977, 
    542, 
    920, 
    1179, 
    529, 
    528, 
    1110, 
    528, 
    980, 
    1110, 
    1110, 
    980, 
    532, 
    530, 
    1110, 
    531, 
    530, 
    529, 
    1110, 
    532, 
    531, 
    1110, 
    980, 
    653, 
    1147, 
    532, 
    980, 
    654, 
    528, 
    653, 
    980, 
    980, 
    1147, 
    654, 
    1147, 
    527, 
    2230, 
    654, 
    1147, 
    533, 
    653, 
    527, 
    1147, 
    1147, 
    2230, 
    533, 
    2230, 
    526, 
    1306, 
    3160, 
    1503, 
    1306, 
    526, 
    3160, 
    1306, 
    1889, 
    1503, 
    3160, 
    4089, 
    3547, 
    1889, 
    524, 
    4089, 
    525, 
    4593, 
    4392, 
    1048, 
    4089, 
    4593, 
    4304, 
    524, 
    523, 
    4593, 
    1373, 
    2035, 
    4904, 
    1503, 
    5077, 
    2297, 
    4494, 
    977, 
    1761, 
    970, 
    5427, 
    1911, 
    2008, 
    977, 
    4494, 
    5427, 
    5130, 
    2008, 
    1911, 
    5427, 
    4494, 
    4986, 
    5130, 
    5427, 
    1754, 
    4986, 
    970, 
    4331, 
    810, 
    5130, 
    544, 
    543, 
    2008, 
    543, 
    542, 
    1179, 
    2230, 
    527, 
    526, 
    534, 
    2230, 
    1306, 
    534, 
    533, 
    2230, 
    2297, 
    1761, 
    836, 
    1306, 
    2297, 
    534, 
    1306, 
    1503, 
    2297, 
    525, 
    1889, 
    3160, 
    1761, 
    977, 
    2214, 
    534, 
    2297, 
    836, 
    1503, 
    1470, 
    5077, 
    4494, 
    5077, 
    1911, 
    526, 
    525, 
    3160, 
    4904, 
    2035, 
    861, 
    1889, 
    4904, 
    1503, 
    1889, 
    3547, 
    4904, 
    861, 
    1671, 
    4598, 
    2607, 
    5714, 
    2996, 
    5070, 
    3032, 
    2645, 
    3967, 
    5070, 
    2672, 
    6346, 
    2889, 
    3234, 
    5070, 
    6346, 
    5352, 
    3967, 
    2889, 
    6346, 
    2696, 
    3967, 
    2672, 
    6346, 
    3234, 
    6090, 
    3017, 
    3350, 
    2472, 
    5352, 
    5257, 
    3364, 
    3967, 
    6346, 
    5070, 
    6090, 
    5257, 
    5352, 
    6346, 
    6090, 
    5352, 
    3234, 
    3545, 
    6090, 
    3654, 
    3234, 
    2889, 
    3350, 
    3654, 
    2889, 
    3178, 
    2996, 
    3654, 
    3665, 
    3936, 
    3586, 
    3894, 
    3625, 
    3042, 
    3375, 
    3894, 
    3042, 
    2453, 
    2871, 
    3894, 
    4234, 
    4521, 
    4962, 
    3221, 
    3319, 
    3625, 
    5351, 
    791, 
    4532, 
    3319, 
    5351, 
    2658, 
    3319, 
    2000, 
    5351, 
    4532, 
    1621, 
    4440, 
    2645, 
    4532, 
    4440, 
    4332, 
    2658, 
    5351, 
    5350, 
    974, 
    1692, 
    2245, 
    5350, 
    1692, 
    2245, 
    4480, 
    5350, 
    4181, 
    2939, 
    2533, 
    4500, 
    3944, 
    4181, 
    1304, 
    4500, 
    4181, 
    1989, 
    4675, 
    4500, 
    3674, 
    3280, 
    3944, 
    4123, 
    3364, 
    3859, 
    3545, 
    3234, 
    2996, 
    3054, 
    4301, 
    4776, 
    4608, 
    6090, 
    3545, 
    5352, 
    3364, 
    3032, 
    4608, 
    5257, 
    6090, 
    5148, 
    3665, 
    5257, 
    5148, 
    3936, 
    3665, 
    3364, 
    5257, 
    3665, 
    4608, 
    5007, 
    5148, 
    5714, 
    4608, 
    3545, 
    2673, 
    3054, 
    4776, 
    3586, 
    3859, 
    3665, 
    3674, 
    3586, 
    3280, 
    3375, 
    3859, 
    3586, 
    3032, 
    5070, 
    5352, 
    2672, 
    5070, 
    2645, 
    4176, 
    2844, 
    2939, 
    3936, 
    4176, 
    3280, 
    5007, 
    4608, 
    4776, 
    3586, 
    3936, 
    3280, 
    5148, 
    5257, 
    4608, 
    4041, 
    3054, 
    2673, 
    4728, 
    4564, 
    2527, 
    5046, 
    4644, 
    4820, 
    5269, 
    5046, 
    4901, 
    5171, 
    5269, 
    4901, 
    4618, 
    4419, 
    5269, 
    5367, 
    4207, 
    5096, 
    5316, 
    3178, 
    2826, 
    4564, 
    5316, 
    2732, 
    4973, 
    5216, 
    5316, 
    4728, 
    4973, 
    4564, 
    4820, 
    5089, 
    5216, 
    4901, 
    4820, 
    4973, 
    5171, 
    4901, 
    4728, 
    5153, 
    5171, 
    4728, 
    4787, 
    4618, 
    5171, 
    5367, 
    4419, 
    4207, 
    6109, 
    5367, 
    5096, 
    5269, 
    4419, 
    5367, 
    4644, 
    4947, 
    5089, 
    4947, 
    4644, 
    4463, 
    2542, 
    4947, 
    4463, 
    4041, 
    2607, 
    5089, 
    4901, 
    4973, 
    4728, 
    5343, 
    3387, 
    3054, 
    2542, 
    5343, 
    4041, 
    2542, 
    4475, 
    5343, 
    4176, 
    2939, 
    3280, 
    3072, 
    3053, 
    1140, 
    2392, 
    4854, 
    1877, 
    2696, 
    3053, 
    3072, 
    2472, 
    3967, 
    2696, 
    2672, 
    4440, 
    3053, 
    3053, 
    2191, 
    1140, 
    1877, 
    3072, 
    1140, 
    2672, 
    2645, 
    4440, 
    4000, 
    2060, 
    1412, 
    1621, 
    4000, 
    2191, 
    1621, 
    4592, 
    4000, 
    4181, 
    2295, 
    1304, 
    4123, 
    4332, 
    3032, 
    4809, 
    2732, 
    2826, 
    4656, 
    4475, 
    2947, 
    3593, 
    4832, 
    3287, 
    3952, 
    3683, 
    4656, 
    4685, 
    3194, 
    2844, 
    4686, 
    4504, 
    4505, 
    3683, 
    4686, 
    4505, 
    3952, 
    1474, 
    4686, 
    2098, 
    974, 
    4504, 
    3054, 
    4041, 
    5343, 
    1759, 
    2295, 
    2533, 
    4592, 
    1621, 
    791, 
    3439, 
    4592, 
    791, 
    911, 
    4000, 
    4592, 
    2191, 
    4000, 
    4300, 
    911, 
    2060, 
    4000, 
    6305, 
    3172, 
    5105, 
    2954, 
    6305, 
    2549, 
    3490, 
    3172, 
    6305, 
    2229, 
    3775, 
    1203, 
    3775, 
    4038, 
    5795, 
    6305, 
    4449, 
    3490, 
    2229, 
    1671, 
    4038, 
    911, 
    5072, 
    5105, 
    5072, 
    1705, 
    3354, 
    1892, 
    1156, 
    2355, 
    2403, 
    1892, 
    1399, 
    5714, 
    2607, 
    2673, 
    4608, 
    5714, 
    2673, 
    3545, 
    2996, 
    5714, 
    3350, 
    2826, 
    3654, 
    4564, 
    2732, 
    4367, 
    5153, 
    4787, 
    5171, 
    4884, 
    5153, 
    2527, 
    2522, 
    4707, 
    5153, 
    4973, 
    5316, 
    4564, 
    3234, 
    3654, 
    2996, 
    2826, 
    2732, 
    5316, 
    3654, 
    2826, 
    3178, 
    2472, 
    3350, 
    2889, 
    3017, 
    4809, 
    3350, 
    5008, 
    3017, 
    2472, 
    2696, 
    5008, 
    2472, 
    4854, 
    2630, 
    5008, 
    2630, 
    4444, 
    4632, 
    4901, 
    5046, 
    4820, 
    4156, 
    4367, 
    2508, 
    5216, 
    4973, 
    4820, 
    5857, 
    5216, 
    5089, 
    2607, 
    5857, 
    5089, 
    2607, 
    2996, 
    5857, 
    3178, 
    5316, 
    5216, 
    4504, 
    974, 
    3194, 
    4854, 
    2392, 
    4369, 
    3017, 
    5008, 
    2630, 
    3072, 
    1877, 
    4854, 
    4444, 
    2920, 
    4632, 
    4369, 
    4444, 
    2630, 
    3262, 
    2920, 
    4444, 
    956, 
    3569, 
    2092, 
    2581, 
    3907, 
    3262, 
    4809, 
    2508, 
    2732, 
    3350, 
    4809, 
    2826, 
    4632, 
    2508, 
    4809, 
    2630, 
    4632, 
    3017, 
    2920, 
    2508, 
    4632, 
    4444, 
    4232, 
    3262, 
    4854, 
    4369, 
    2630, 
    1460, 
    4232, 
    4369, 
    4541, 
    2692, 
    3579, 
    4709, 
    4541, 
    3273, 
    3277, 
    3583, 
    4541, 
    4367, 
    4156, 
    2935, 
    2527, 
    4367, 
    2935, 
    2732, 
    2508, 
    4367, 
    3583, 
    2692, 
    4541, 
    4156, 
    3907, 
    3277, 
    3622, 
    3315, 
    2492, 
    2581, 
    3622, 
    3583, 
    2581, 
    2974, 
    3622, 
    3569, 
    2581, 
    3262, 
    1742, 
    2974, 
    956, 
    1742, 
    2284, 
    3315, 
    2974, 
    3315, 
    3622, 
    2092, 
    3569, 
    4232, 
    4300, 
    1877, 
    1140, 
    2392, 
    1188, 
    1460, 
    4505, 
    4685, 
    4301, 
    4039, 
    3778, 
    2772, 
    2203, 
    4039, 
    1640, 
    2203, 
    1158, 
    4117, 
    4903, 
    4556, 
    2011, 
    2321, 
    5213, 
    1335, 
    1692, 
    892, 
    4903, 
    892, 
    2050, 
    4556, 
    1474, 
    2403, 
    2050, 
    5008, 
    2696, 
    3072, 
    2889, 
    3967, 
    2472, 
    2672, 
    3053, 
    2696, 
    2403, 
    1399, 
    2050, 
    4848, 
    1008, 
    3514, 
    5123, 
    4848, 
    1229, 
    1784, 
    1008, 
    4848, 
    2245, 
    5123, 
    1229, 
    4480, 
    2245, 
    1229, 
    2980, 
    4480, 
    1229, 
    1759, 
    5350, 
    4480, 
    5213, 
    4903, 
    1335, 
    5123, 
    5213, 
    2321, 
    1692, 
    4903, 
    5213, 
    5920, 
    2435, 
    2855, 
    2652, 
    5740, 
    2432, 
    2652, 
    5401, 
    5740, 
    2653, 
    4990, 
    2432, 
    5431, 
    790, 
    1620, 
    5123, 
    2321, 
    1784, 
    4848, 
    5123, 
    1784, 
    2245, 
    5213, 
    5123, 
    3455, 
    2011, 
    2715, 
    2245, 
    1692, 
    5213, 
    2307, 
    2632, 
    3743, 
    2307, 
    1317, 
    2632, 
    3940, 
    3670, 
    2431, 
    3200, 
    4178, 
    2851, 
    3515, 
    3670, 
    3940, 
    3671, 
    3131, 
    3370, 
    3795, 
    3941, 
    3515, 
    3455, 
    3131, 
    3671, 
    2768, 
    3370, 
    3131, 
    2768, 
    3038, 
    3370, 
    3940, 
    2431, 
    2851, 
    2852, 
    5920, 
    3201, 
    3201, 
    5920, 
    3670, 
    5326, 
    773, 
    1989, 
    1508, 
    1540, 
    688, 
    2421, 
    1915, 
    2134, 
    1540, 
    2421, 
    2134, 
    3002, 
    2114, 
    3200, 
    2114, 
    1508, 
    688, 
    1939, 
    3514, 
    688, 
    4473, 
    2564, 
    3025, 
    4763, 
    4389, 
    1999, 
    5968, 
    4934, 
    4763, 
    5431, 
    5968, 
    4763, 
    5347, 
    4473, 
    6444, 
    4473, 
    5347, 
    4214, 
    4473, 
    5133, 
    5625, 
    4934, 
    4389, 
    4763, 
    4934, 
    4589, 
    4389, 
    3723, 
    3433, 
    5133, 
    4236, 
    5248, 
    4447, 
    5827, 
    4933, 
    5071, 
    5248, 
    5827, 
    5132, 
    5248, 
    6005, 
    5827, 
    4447, 
    5248, 
    5132, 
    6005, 
    4761, 
    4933, 
    5142, 
    6005, 
    5248, 
    5142, 
    5868, 
    6005, 
    1620, 
    2190, 
    4214, 
    4178, 
    1008, 
    1784, 
    3515, 
    3671, 
    3201, 
    2411, 
    571, 
    570, 
    6639, 
    3577, 
    564, 
    1489, 
    2519, 
    2411, 
    2682, 
    1445, 
    2384, 
    4690, 
    2682, 
    2384, 
    1369, 
    855, 
    2682, 
    2682, 
    855, 
    2081, 
    2027, 
    2284, 
    846, 
    2951, 
    3291, 
    2907, 
    757, 
    4847, 
    1979, 
    4924, 
    4750, 
    4674, 
    757, 
    5061, 
    4847, 
    5778, 
    4750, 
    4924, 
    5061, 
    5778, 
    4924, 
    3639, 
    3909, 
    5872, 
    3622, 
    2492, 
    2692, 
    1742, 
    3315, 
    2974, 
    2284, 
    2907, 
    3315, 
    4556, 
    815, 
    2011, 
    1335, 
    4903, 
    2011, 
    2050, 
    3459, 
    4556, 
    1474, 
    2050, 
    892, 
    1399, 
    3459, 
    2050, 
    2098, 
    1474, 
    892, 
    1692, 
    2098, 
    892, 
    3194, 
    1759, 
    2533, 
    4023, 
    1077, 
    3187, 
    2837, 
    4023, 
    3187, 
    3758, 
    4237, 
    4448, 
    1156, 
    1832, 
    2355, 
    1156, 
    2201, 
    1832, 
    1566, 
    2154, 
    811, 
    2009, 
    1566, 
    811, 
    4832, 
    1892, 
    2403, 
    4656, 
    4832, 
    3952, 
    4656, 
    3287, 
    4832, 
    1333, 
    727, 
    2009, 
    727, 
    4286, 
    5019, 
    3459, 
    815, 
    4556, 
    3459, 
    4237, 
    1640, 
    1892, 
    2355, 
    1399, 
    4448, 
    4023, 
    3758, 
    2355, 
    4448, 
    4237, 
    1832, 
    4023, 
    4448, 
    4548, 
    4724, 
    5194, 
    3459, 
    2355, 
    4237, 
    815, 
    3459, 
    1640, 
    1399, 
    2355, 
    3459, 
    4277, 
    2496, 
    3511, 
    3741, 
    2410, 
    2962, 
    5127, 
    5242, 
    3452, 
    1901, 
    2410, 
    3741, 
    4034, 
    2496, 
    2808, 
    5127, 
    4034, 
    2808, 
    2618, 
    3005, 
    4258, 
    3712, 
    3882, 
    3417, 
    6185, 
    3612, 
    2653, 
    3038, 
    6185, 
    2653, 
    3882, 
    3612, 
    6185, 
    3417, 
    3882, 
    2768, 
    3712, 
    3612, 
    3882, 
    4011, 
    3712, 
    3417, 
    5642, 
    2823, 
    4206, 
    3712, 
    5642, 
    3978, 
    3175, 
    2823, 
    5642, 
    3306, 
    4634, 
    3612, 
    4272, 
    3835, 
    4648, 
    4648, 
    3835, 
    3561, 
    3916, 
    4272, 
    3646, 
    3916, 
    4048, 
    4272, 
    5199, 
    2100, 
    978, 
    5131, 
    5199, 
    3805, 
    4101, 
    2100, 
    5199, 
    4272, 
    4101, 
    3835, 
    1477, 
    2100, 
    4101, 
    3526, 
    3210, 
    3214, 
    2837, 
    2404, 
    1893, 
    1158, 
    3758, 
    1893, 
    5019, 
    1566, 
    727, 
    4869, 
    4561, 
    4364, 
    2100, 
    4869, 
    4067, 
    1477, 
    4561, 
    4869, 
    3187, 
    2154, 
    4364, 
    3758, 
    4023, 
    2837, 
    2154, 
    1566, 
    4364, 
    4561, 
    2837, 
    3187, 
    5019, 
    4869, 
    4364, 
    1566, 
    5019, 
    4364, 
    4286, 
    4067, 
    5019, 
    2404, 
    2837, 
    4561, 
    5514, 
    3910, 
    3640, 
    2860, 
    5286, 
    3210, 
    4159, 
    3910, 
    5189, 
    1990, 
    4159, 
    1307, 
    3519, 
    3910, 
    4159, 
    2963, 
    5135, 
    5250, 
    4063, 
    2445, 
    3802, 
    5514, 
    6044, 
    3802, 
    2998, 
    2610, 
    5497, 
    4277, 
    4051, 
    2808, 
    2496, 
    4277, 
    2808, 
    3511, 
    3791, 
    4277, 
    2860, 
    1762, 
    2298, 
    1307, 
    4159, 
    5286, 
    3252, 
    2910, 
    4258, 
    5131, 
    3805, 
    3526, 
    3214, 
    5395, 
    3526, 
    3835, 
    4101, 
    5199, 
    5468, 
    2846, 
    2910, 
    5395, 
    5468, 
    3252, 
    3214, 
    3523, 
    5832, 
    3561, 
    5395, 
    3252, 
    978, 
    3805, 
    5199, 
    3805, 
    2860, 
    3526, 
    3561, 
    3835, 
    5131, 
    978, 
    1762, 
    3805, 
    6044, 
    3334, 
    2998, 
    5497, 
    6044, 
    2998, 
    4063, 
    3802, 
    6044, 
    2846, 
    5832, 
    2445, 
    5514, 
    3640, 
    3334, 
    3523, 
    5514, 
    3802, 
    3523, 
    5189, 
    5514, 
    3210, 
    3523, 
    3214, 
    5348, 
    3519, 
    3610, 
    5514, 
    5189, 
    3910, 
    5189, 
    3210, 
    5286, 
    4565, 
    4370, 
    4981, 
    1581, 
    4565, 
    747, 
    4391, 
    4370, 
    4565, 
    2166, 
    4391, 
    1581, 
    2664, 
    4370, 
    4391, 
    5121, 
    1669, 
    4495, 
    4391, 
    4565, 
    1581, 
    1363, 
    1974, 
    1275, 
    1363, 
    2027, 
    1974, 
    2337, 
    1979, 
    1363, 
    1799, 
    2337, 
    1275, 
    757, 
    1979, 
    2337, 
    1287, 
    2027, 
    1363, 
    4181, 
    2533, 
    2295, 
    1989, 
    4500, 
    1304, 
    3944, 
    2939, 
    4181, 
    3944, 
    3280, 
    2939, 
    4359, 
    4146, 
    3674, 
    4500, 
    4359, 
    3944, 
    4675, 
    773, 
    4445, 
    3375, 
    3586, 
    3674, 
    3894, 
    3375, 
    4146, 
    3859, 
    3364, 
    3665, 
    3042, 
    3859, 
    3375, 
    3042, 
    4123, 
    3859, 
    2871, 
    3625, 
    3894, 
    4123, 
    3032, 
    3364, 
    2658, 
    4123, 
    3042, 
    2658, 
    4332, 
    4123, 
    2844, 
    2533, 
    2939, 
    4853, 
    4301, 
    4685, 
    4176, 
    4853, 
    2844, 
    4776, 
    4301, 
    4853, 
    5007, 
    4776, 
    4853, 
    3936, 
    5007, 
    4176, 
    3936, 
    5148, 
    5007, 
    4608, 
    2673, 
    4776, 
    2607, 
    4041, 
    2673, 
    2542, 
    2947, 
    4475, 
    3194, 
    2533, 
    2844, 
    4505, 
    3387, 
    3683, 
    4176, 
    5007, 
    4853, 
    3054, 
    3387, 
    4301, 
    974, 
    1759, 
    3194, 
    3474, 
    2778, 
    3138, 
    3593, 
    3474, 
    1156, 
    1892, 
    3593, 
    1156, 
    3287, 
    3762, 
    3593, 
    3593, 
    3762, 
    3474, 
    4832, 
    2403, 
    3952, 
    3762, 
    2778, 
    3474, 
    2947, 
    4027, 
    3287, 
    5451, 
    5375, 
    3117, 
    3287, 
    4027, 
    3762, 
    2947, 
    2542, 
    4253, 
    2098, 
    4686, 
    1474, 
    5375, 
    5278, 
    2751, 
    2947, 
    4253, 
    4027, 
    2542, 
    4041, 
    4947, 
    3583, 
    3622, 
    2692, 
    1637, 
    1077, 
    2201, 
    2154, 
    1637, 
    811, 
    1077, 
    1832, 
    2201, 
    4237, 
    3758, 
    2203, 
    1640, 
    4237, 
    2203, 
    2355, 
    1832, 
    4448, 
    1754, 
    1920, 
    1664, 
    2220, 
    956, 
    2092, 
    2166, 
    1660, 
    2220, 
    2343, 
    3949, 
    1373, 
    3924, 
    2366, 
    1412, 
    3652, 
    3924, 
    2819, 
    3652, 
    6180, 
    4082, 
    6190, 
    6180, 
    3349, 
    4082, 
    3817, 
    1845, 
    3652, 
    4082, 
    3924, 
    3540, 
    3817, 
    4082, 
    3172, 
    3652, 
    2819, 
    1581, 
    1660, 
    2166, 
    1581, 
    846, 
    1660, 
    5936, 
    2000, 
    1318, 
    911, 
    4592, 
    1705, 
    791, 
    2000, 
    3439, 
    3674, 
    4146, 
    3375, 
    5159, 
    2181, 
    1124, 
    4234, 
    2710, 
    4521, 
    4146, 
    6256, 
    2453, 
    4146, 
    4359, 
    6256, 
    1608, 
    2181, 
    2710, 
    5150, 
    1242, 
    2256, 
    2308, 
    5150, 
    1318, 
    2308, 
    4309, 
    5150, 
    5915, 
    1772, 
    990, 
    1949, 
    5915, 
    4050, 
    4309, 
    1772, 
    5915, 
    5150, 
    4309, 
    1242, 
    2308, 
    1772, 
    4309, 
    3221, 
    2308, 
    1318, 
    2000, 
    3319, 
    1318, 
    2871, 
    5101, 
    5227, 
    5227, 
    5101, 
    4110, 
    3221, 
    5227, 
    2308, 
    3221, 
    2871, 
    5227, 
    4309, 
    5915, 
    1949, 
    4962, 
    2871, 
    2453, 
    5227, 
    4110, 
    1772, 
    4962, 
    5101, 
    2871, 
    4324, 
    4110, 
    5101, 
    4962, 
    4324, 
    5101, 
    4234, 
    4962, 
    2453, 
    4521, 
    4324, 
    4962, 
    2181, 
    5159, 
    2710, 
    5159, 
    4524, 
    6116, 
    2710, 
    5159, 
    4521, 
    1124, 
    4524, 
    5159, 
    1124, 
    1867, 
    4524, 
    990, 
    1772, 
    4110, 
    5415, 
    2134, 
    3930, 
    5326, 
    5415, 
    773, 
    1540, 
    2134, 
    5415, 
    1772, 
    2308, 
    5227, 
    3930, 
    2181, 
    1608, 
    4578, 
    1124, 
    2181, 
    3930, 
    4578, 
    2181, 
    1042, 
    1197, 
    4578, 
    1949, 
    1242, 
    4309, 
    990, 
    4050, 
    5915, 
    707, 
    2325, 
    5087, 
    1986, 
    767, 
    3852, 
    1514, 
    1986, 
    851, 
    1514, 
    2635, 
    6020, 
    6494, 
    2256, 
    1242, 
    4526, 
    6020, 
    6494, 
    2635, 
    3354, 
    3657, 
    2426, 
    4590, 
    1514, 
    3354, 
    1705, 
    3657, 
    4592, 
    3439, 
    1705, 
    1986, 
    1514, 
    6020, 
    3439, 
    2256, 
    1705, 
    3439, 
    5936, 
    2256, 
    4526, 
    1604, 
    767, 
    1581, 
    747, 
    846, 
    4501, 
    3949, 
    2343, 
    2659, 
    4501, 
    1809, 
    2659, 
    3043, 
    4501, 
    3678, 
    3376, 
    3380, 
    5598, 
    4392, 
    522, 
    1546, 
    5598, 
    521, 
    1546, 
    2138, 
    5598, 
    4593, 
    1048, 
    1809, 
    522, 
    4392, 
    523, 
    2138, 
    1048, 
    4392, 
    522, 
    521, 
    5598, 
    5944, 
    6106, 
    2608, 
    5809, 
    5554, 
    5656, 
    6451, 
    6068, 
    5944, 
    6422, 
    6451, 
    5656, 
    6517, 
    5001, 
    6068, 
    6422, 
    6517, 
    6451, 
    6422, 
    5531, 
    6517, 
    3331, 
    2994, 
    5809, 
    5001, 
    520, 
    3825, 
    520, 
    1546, 
    521, 
    520, 
    994, 
    3825, 
    2138, 
    4392, 
    5598, 
    516, 
    1322, 
    2311, 
    994, 
    519, 
    518, 
    517, 
    994, 
    518, 
    1669, 
    859, 
    4040, 
    6683, 
    509, 
    508, 
    6683, 
    510, 
    509, 
    507, 
    6684, 
    508, 
    6684, 
    510, 
    6683, 
    6646, 
    6684, 
    507, 
    1930, 
    6646, 
    507, 
    6684, 
    6683, 
    508, 
    511, 
    6684, 
    6646, 
    511, 
    510, 
    6684, 
    1388, 
    1930, 
    506, 
    6602, 
    512, 
    669, 
    513, 
    6602, 
    514, 
    513, 
    512, 
    6602, 
    512, 
    511, 
    669, 
    1930, 
    511, 
    6646, 
    506, 
    1930, 
    507, 
    1388, 
    2195, 
    2316, 
    6694, 
    505, 
    651, 
    687, 
    6694, 
    651, 
    652, 
    505, 
    6694, 
    687, 
    651, 
    504, 
    6694, 
    687, 
    4623, 
    687, 
    876, 
    4623, 
    503, 
    1464, 
    504, 
    4887, 
    2638, 
    3024, 
    1464, 
    4219, 
    876, 
    4797, 
    1512, 
    2424, 
    5398, 
    4797, 
    4219, 
    1464, 
    5398, 
    4219, 
    3198, 
    2849, 
    5398, 
    2849, 
    1512, 
    4797, 
    669, 
    514, 
    6602, 
    652, 
    6694, 
    4623, 
    6230, 
    2117, 
    2849, 
    4623, 
    876, 
    960, 
    1388, 
    4623, 
    960, 
    506, 
    652, 
    4623, 
    687, 
    504, 
    1464, 
    3552, 
    669, 
    2316, 
    2003, 
    6211, 
    796, 
    514, 
    669, 
    3552, 
    4306, 
    1669, 
    4040, 
    1625, 
    3731, 
    4306, 
    2933, 
    2525, 
    2646, 
    4177, 
    2933, 
    2646, 
    4287, 
    4495, 
    2646, 
    2227, 
    1201, 
    4177, 
    1201, 
    1918, 
    2933, 
    1536, 
    946, 
    2085, 
    5528, 
    3588, 
    3860, 
    5014, 
    6421, 
    678, 
    1426, 
    2532, 
    5743, 
    4294, 
    946, 
    1536, 
    1106, 
    4294, 
    1536, 
    1106, 
    6227, 
    4294, 
    4294, 
    1034, 
    1732, 
    1979, 
    1287, 
    1363, 
    1275, 
    2337, 
    1363, 
    5517, 
    5061, 
    1593, 
    3333, 
    5517, 
    2997, 
    3333, 
    5778, 
    5517, 
    1799, 
    1593, 
    757, 
    2278, 
    1799, 
    1275, 
    3365, 
    3806, 
    4068, 
    1974, 
    3215, 
    1275, 
    5972, 
    747, 
    4565, 
    1732, 
    1034, 
    2278, 
    1034, 
    1593, 
    1799, 
    1930, 
    669, 
    511, 
    4623, 
    1388, 
    506, 
    960, 
    2195, 
    1388, 
    4040, 
    859, 
    1322, 
    2003, 
    4040, 
    1322, 
    2003, 
    4306, 
    4040, 
    5814, 
    6231, 
    5122, 
    6068, 
    5001, 
    3825, 
    1371, 
    6106, 
    3825, 
    5944, 
    5809, 
    6451, 
    859, 
    1669, 
    5121, 
    4495, 
    4177, 
    2646, 
    4287, 
    3033, 
    4068, 
    1201, 
    2933, 
    4177, 
    2525, 
    3033, 
    2646, 
    3215, 
    3527, 
    3937, 
    4068, 
    3033, 
    3365, 
    2994, 
    4068, 
    2605, 
    2994, 
    4287, 
    4068, 
    5003, 
    4800, 
    3815, 
    2879, 
    5003, 
    2461, 
    4954, 
    4800, 
    5003, 
    946, 
    5094, 
    2879, 
    3582, 
    3854, 
    4954, 
    3666, 
    3582, 
    3276, 
    3365, 
    3033, 
    3854, 
    6211, 
    2858, 
    514, 
    796, 
    6211, 
    3552, 
    2003, 
    2858, 
    6211, 
    4306, 
    2003, 
    796, 
    2858, 
    515, 
    514, 
    1322, 
    2858, 
    2003, 
    1322, 
    515, 
    2858, 
    1500, 
    476, 
    1162, 
    1500, 
    478, 
    477, 
    476, 
    1500, 
    477, 
    6302, 
    4921, 
    2074, 
    1162, 
    6302, 
    1500, 
    1162, 
    1644, 
    6302, 
    500, 
    499, 
    6606, 
    6605, 
    499, 
    498, 
    6609, 
    6605, 
    498, 
    5163, 
    6609, 
    498, 
    502, 
    6605, 
    6609, 
    6606, 
    499, 
    6605, 
    501, 
    6606, 
    6605, 
    501, 
    500, 
    6606, 
    501, 
    6605, 
    502, 
    5163, 
    502, 
    6609, 
    5163, 
    497, 
    2486, 
    6700, 
    495, 
    2486, 
    496, 
    6700, 
    497, 
    496, 
    495, 
    6700, 
    497, 
    6700, 
    2486, 
    1770, 
    494, 
    493, 
    6669, 
    491, 
    2306, 
    492, 
    6669, 
    493, 
    492, 
    491, 
    6669, 
    491, 
    1814, 
    2306, 
    6610, 
    488, 
    487, 
    6610, 
    489, 
    488, 
    6611, 
    6610, 
    487, 
    1814, 
    6611, 
    487, 
    490, 
    6610, 
    6611, 
    490, 
    489, 
    6610, 
    1814, 
    490, 
    6611, 
    6586, 
    486, 
    485, 
    484, 
    6586, 
    485, 
    484, 
    1138, 
    6649, 
    486, 
    6586, 
    6649, 
    1814, 
    6649, 
    1138, 
    480, 
    6670, 
    481, 
    6671, 
    479, 
    667, 
    6670, 
    6671, 
    482, 
    6670, 
    480, 
    6671, 
    481, 
    6670, 
    482, 
    480, 
    479, 
    6671, 
    650, 
    6671, 
    667, 
    650, 
    667, 
    1527, 
    6671, 
    650, 
    482, 
    1500, 
    479, 
    478, 
    1992, 
    1162, 
    476, 
    3150, 
    2905, 
    1992, 
    475, 
    3150, 
    476, 
    1561, 
    2905, 
    3150, 
    779, 
    1644, 
    1992, 
    1644, 
    818, 
    2406, 
    1992, 
    1644, 
    1162, 
    779, 
    818, 
    1644, 
    5880, 
    5173, 
    779, 
    721, 
    5880, 
    2905, 
    1394, 
    5173, 
    5880, 
    6156, 
    4544, 
    4711, 
    3830, 
    6156, 
    721, 
    6282, 
    2556, 
    4544, 
    3830, 
    6282, 
    6156, 
    3830, 
    3557, 
    6282, 
    1253, 
    4888, 
    5173, 
    4888, 
    885, 
    4006, 
    3995, 
    4133, 
    3297, 
    3122, 
    1103, 
    1852, 
    3122, 
    2755, 
    3246, 
    2372, 
    3297, 
    1852, 
    3297, 
    4133, 
    3122, 
    3830, 
    721, 
    1561, 
    2755, 
    6282, 
    3557, 
    6282, 
    4544, 
    6156, 
    4133, 
    2556, 
    2755, 
    3122, 
    4133, 
    2755, 
    6074, 
    3275, 
    3581, 
    3995, 
    4223, 
    4133, 
    3995, 
    2501, 
    4223, 
    4095, 
    5169, 
    2501, 
    6466, 
    3853, 
    5816, 
    4711, 
    6466, 
    5816, 
    5739, 
    3581, 
    6466, 
    5169, 
    3581, 
    3275, 
    2501, 
    5169, 
    3275, 
    3829, 
    3556, 
    6052, 
    6169, 
    3245, 
    2904, 
    3853, 
    6169, 
    4119, 
    6052, 
    3245, 
    6169, 
    3830, 
    1561, 
    4022, 
    6230, 
    1012, 
    2117, 
    4938, 
    4769, 
    6230, 
    981, 
    4938, 
    1602, 
    981, 
    5255, 
    4938, 
    1786, 
    1012, 
    4769, 
    5255, 
    1786, 
    4769, 
    4735, 
    5255, 
    981, 
    2323, 
    1786, 
    5255, 
    2102, 
    4735, 
    981, 
    3499, 
    1130, 
    1870, 
    1339, 
    2629, 
    5429, 
    1339, 
    2013, 
    2629, 
    3499, 
    2629, 
    1130, 
    4006, 
    1130, 
    2185, 
    1690, 
    4006, 
    885, 
    1690, 
    3016, 
    4006, 
    1253, 
    5816, 
    6075, 
    3016, 
    1870, 
    1130, 
    923, 
    3016, 
    1690, 
    923, 
    1222, 
    3016, 
    2085, 
    678, 
    1536, 
    4600, 
    1870, 
    2388, 
    3685, 
    6279, 
    4600, 
    4045, 
    3785, 
    3388, 
    3502, 
    1012, 
    3954, 
    5429, 
    2323, 
    1339, 
    3499, 
    5429, 
    2629, 
    3782, 
    2323, 
    5429, 
    6279, 
    3782, 
    3499, 
    4600, 
    6279, 
    3499, 
    3685, 
    3954, 
    6279, 
    1786, 
    2323, 
    3782, 
    2388, 
    1222, 
    5014, 
    3016, 
    1222, 
    1870, 
    5569, 
    2489, 
    2532, 
    1222, 
    5569, 
    2532, 
    923, 
    4329, 
    6430, 
    1862, 
    2380, 
    1480, 
    4888, 
    4006, 
    2185, 
    1770, 
    495, 
    494, 
    6669, 
    1770, 
    493, 
    6072, 
    981, 
    1602, 
    1770, 
    6072, 
    2486, 
    1116, 
    981, 
    6072, 
    2013, 
    5317, 
    2629, 
    779, 
    1613, 
    818, 
    779, 
    2905, 
    5880, 
    2486, 
    495, 
    1770, 
    1116, 
    6072, 
    1770, 
    1602, 
    766, 
    5163, 
    5255, 
    4769, 
    4938, 
    5163, 
    498, 
    497, 
    1602, 
    5163, 
    2486, 
    766, 
    503, 
    5163, 
    1527, 
    1138, 
    484, 
    2306, 
    1116, 
    1770, 
    2380, 
    1862, 
    1316, 
    4187, 
    2380, 
    1316, 
    1436, 
    2406, 
    2380, 
    1480, 
    2102, 
    1862, 
    2406, 
    1480, 
    2380, 
    2074, 
    4748, 
    1436, 
    818, 
    2013, 
    2406, 
    4735, 
    2323, 
    5255, 
    2306, 
    1770, 
    6669, 
    1862, 
    2306, 
    1316, 
    1862, 
    1116, 
    2306, 
    1527, 
    483, 
    650, 
    4921, 
    4748, 
    2074, 
    1644, 
    4921, 
    6302, 
    1644, 
    2406, 
    4921, 
    1814, 
    491, 
    490, 
    6649, 
    1814, 
    487, 
    486, 
    6649, 
    487, 
    6586, 
    484, 
    6649, 
    1138, 
    1316, 
    1814, 
    1814, 
    1316, 
    2306, 
    1527, 
    1436, 
    4187, 
    483, 
    1527, 
    484, 
    667, 
    2074, 
    1527, 
    5317, 
    818, 
    1613, 
    4735, 
    2013, 
    1339, 
    1480, 
    2406, 
    2013, 
    4187, 
    1436, 
    2380, 
    1138, 
    4187, 
    1316, 
    1138, 
    1527, 
    4187, 
    6302, 
    479, 
    1500, 
    1527, 
    2074, 
    1436, 
    667, 
    479, 
    2074, 
    6072, 
    1602, 
    2486, 
    5880, 
    721, 
    1394, 
    476, 
    3150, 
    1992, 
    1561, 
    721, 
    2905, 
    4045, 
    1450, 
    2085, 
    1222, 
    2388, 
    1870, 
    1222, 
    1426, 
    5014, 
    502, 
    5163, 
    503, 
    4748, 
    2406, 
    1436, 
    479, 
    6302, 
    2074, 
    4921, 
    2406, 
    4748, 
    1599, 
    6220, 
    763, 
    1322, 
    516, 
    515, 
    514, 
    3552, 
    6211, 
    859, 
    2033, 
    1322, 
    1589, 
    474, 
    473, 
    3150, 
    1070, 
    1561, 
    3150, 
    475, 
    1070, 
    475, 
    474, 
    1070, 
    5080, 
    466, 
    1283, 
    4904, 
    861, 
    1470, 
    1503, 
    4904, 
    1470, 
    4501, 
    2343, 
    1809, 
    4680, 
    3949, 
    4501, 
    3678, 
    3973, 
    4203, 
    3376, 
    3678, 
    4680, 
    3380, 
    3708, 
    3678, 
    4304, 
    1809, 
    2343, 
    4089, 
    4304, 
    3547, 
    4089, 
    524, 
    4593, 
    2166, 
    2706, 
    4391, 
    523, 
    4392, 
    4593, 
    3825, 
    994, 
    1371, 
    4287, 
    2994, 
    3331, 
    5121, 
    4287, 
    3331, 
    5121, 
    4495, 
    4287, 
    2608, 
    5121, 
    3331, 
    2608, 
    859, 
    5121, 
    1669, 
    2227, 
    4495, 
    2646, 
    3033, 
    4287, 
    520, 
    5001, 
    1546, 
    1371, 
    517, 
    2311, 
    6170, 
    2659, 
    1048, 
    5944, 
    3331, 
    5809, 
    3043, 
    2659, 
    5531, 
    994, 
    517, 
    1371, 
    2608, 
    6106, 
    2033, 
    859, 
    2608, 
    2033, 
    5809, 
    2994, 
    5554, 
    519, 
    994, 
    520, 
    2311, 
    1322, 
    2033, 
    1371, 
    2311, 
    2033, 
    517, 
    516, 
    2311, 
    1464, 
    876, 
    687, 
    6230, 
    4769, 
    1012, 
    3198, 
    6230, 
    2849, 
    6401, 
    766, 
    4938, 
    3198, 
    6401, 
    6230, 
    3198, 
    503, 
    6401, 
    2849, 
    2117, 
    1512, 
    503, 
    3198, 
    1464, 
    4938, 
    766, 
    1602, 
    4797, 
    5398, 
    2849, 
    503, 
    766, 
    6401, 
    4797, 
    2424, 
    2638, 
    4887, 
    4797, 
    2638, 
    3854, 
    4800, 
    4954, 
    2933, 
    4437, 
    2525, 
    4659, 
    3785, 
    2461, 
    4079, 
    4835, 
    3815, 
    3502, 
    3785, 
    4659, 
    1012, 
    3502, 
    2117, 
    4659, 
    2461, 
    3815, 
    3685, 
    3785, 
    3502, 
    3685, 
    3388, 
    3785, 
    3954, 
    3782, 
    6279, 
    3502, 
    3954, 
    3685, 
    1012, 
    1786, 
    3954, 
    2388, 
    1450, 
    3388, 
    4045, 
    2085, 
    2879, 
    1464, 
    3198, 
    5398, 
    4835, 
    4659, 
    3815, 
    1918, 
    1201, 
    3024, 
    2316, 
    669, 
    1930, 
    1388, 
    2316, 
    1930, 
    1625, 
    796, 
    3552, 
    1106, 
    2997, 
    6227, 
    5014, 
    1426, 
    6421, 
    1450, 
    5014, 
    678, 
    1450, 
    2388, 
    5014, 
    4042, 
    4268, 
    2869, 
    3114, 
    3730, 
    3994, 
    4794, 
    1005, 
    2609, 
    1557, 
    3929, 
    4540, 
    3443, 
    1822, 
    2352, 
    3730, 
    3443, 
    2352, 
    3868, 
    4259, 
    4467, 
    3730, 
    3114, 
    3443, 
    1391, 
    3730, 
    2352, 
    1391, 
    2044, 
    4944, 
    2747, 
    2752, 
    4885, 
    2969, 
    2574, 
    2752, 
    3869, 
    3096, 
    3600, 
    4140, 
    3869, 
    3600, 
    3885, 
    4132, 
    3869, 
    3982, 
    4626, 
    6174, 
    4953, 
    2894, 
    2702, 
    3424, 
    4953, 
    3096, 
    4799, 
    2478, 
    4953, 
    2955, 
    3294, 
    2969, 
    5914, 
    5543, 
    5721, 
    6417, 
    6544, 
    6461, 
    6134, 
    6276, 
    6339, 
    6539, 
    6355, 
    6476, 
    6540, 
    6365, 
    6539, 
    6417, 
    6461, 
    6366, 
    6417, 
    6468, 
    6544, 
    5914, 
    6417, 
    6366, 
    5780, 
    5618, 
    6468, 
    6482, 
    6355, 
    6539, 
    6460, 
    6482, 
    6365, 
    5695, 
    5841, 
    6482, 
    6377, 
    6442, 
    6328, 
    6200, 
    5644, 
    5800, 
    5914, 
    6200, 
    5543, 
    6040, 
    6158, 
    6200, 
    3724, 
    5999, 
    6134, 
    3724, 
    3988, 
    5999, 
    6549, 
    5750, 
    5583, 
    5695, 
    6482, 
    6460, 
    6468, 
    5583, 
    5750, 
    6468, 
    5618, 
    5583, 
    6544, 
    6468, 
    5750, 
    5509, 
    6544, 
    5750, 
    6460, 
    6461, 
    6544, 
    6417, 
    5780, 
    6468, 
    5934, 
    5721, 
    5543, 
    5505, 
    5618, 
    5780, 
    5505, 
    2955, 
    5618, 
    5538, 
    3435, 
    4804, 
    5538, 
    3724, 
    3435, 
    4441, 
    5538, 
    2733, 
    4441, 
    3988, 
    5538, 
    5495, 
    3988, 
    4441, 
    5004, 
    5495, 
    4227, 
    4215, 
    3988, 
    5495, 
    1955, 
    5147, 
    4001, 
    5828, 
    6046, 
    3868, 
    5492, 
    6303, 
    5682, 
    4429, 
    4622, 
    5788, 
    6303, 
    4429, 
    5788, 
    5999, 
    5492, 
    5644, 
    6237, 
    6158, 
    6276, 
    5644, 
    6237, 
    5999, 
    6200, 
    6158, 
    6237, 
    4958, 
    3432, 
    3103, 
    2736, 
    4958, 
    3106, 
    2736, 
    3818, 
    5098, 
    5172, 
    1822, 
    3443, 
    930, 
    2112, 
    1504, 
    3729, 
    4400, 
    2319, 
    4768, 
    3479, 
    3765, 
    4599, 
    4768, 
    3765, 
    3113, 
    2746, 
    4937, 
    2512, 
    6096, 
    6391, 
    3442, 
    4768, 
    4599, 
    4147, 
    4239, 
    3897, 
    3729, 
    4599, 
    4400, 
    3159, 
    5318, 
    3479, 
    4400, 
    2609, 
    1782, 
    3442, 
    4599, 
    3729, 
    4032, 
    2609, 
    4400, 
    5090, 
    4032, 
    3765, 
    5090, 
    4949, 
    4032, 
    5983, 
    6492, 
    4949, 
    6492, 
    2771, 
    4794, 
    4949, 
    6492, 
    4794, 
    5983, 
    3458, 
    6492, 
    4794, 
    2771, 
    2112, 
    4032, 
    4949, 
    2609, 
    2609, 
    4949, 
    4794, 
    6492, 
    3458, 
    2771, 
    5806, 
    5983, 
    4949, 
    5806, 
    5940, 
    5983, 
    5829, 
    5518, 
    5683, 
    5573, 
    5705, 
    5483, 
    5573, 
    5536, 
    5705, 
    5940, 
    5806, 
    6014, 
    3747, 
    5940, 
    4010, 
    3747, 
    3458, 
    5983, 
    5219, 
    5318, 
    5715, 
    3765, 
    5219, 
    5090, 
    3159, 
    2804, 
    6391, 
    4872, 
    4147, 
    3897, 
    3580, 
    4872, 
    3274, 
    4701, 
    4147, 
    4872, 
    4529, 
    4360, 
    4701, 
    2952, 
    4529, 
    3292, 
    2528, 
    4557, 
    4529, 
    3747, 
    4010, 
    4360, 
    5022, 
    3897, 
    3629, 
    4701, 
    4360, 
    4147, 
    3292, 
    4701, 
    3580, 
    3292, 
    4529, 
    4701, 
    4010, 
    4239, 
    4147, 
    6232, 
    5536, 
    5573, 
    3747, 
    5983, 
    5940, 
    5090, 
    5219, 
    6014, 
    4949, 
    5090, 
    5806, 
    3765, 
    3479, 
    5219, 
    6096, 
    2512, 
    5493, 
    5683, 
    6096, 
    5493, 
    6391, 
    5318, 
    3159, 
    5518, 
    6391, 
    6096, 
    5518, 
    6513, 
    6391, 
    6513, 
    5318, 
    6391, 
    6513, 
    5715, 
    5318, 
    5705, 
    6513, 
    5518, 
    5705, 
    5536, 
    6513, 
    5536, 
    5940, 
    6014, 
    5219, 
    3479, 
    5318, 
    3629, 
    4955, 
    5022, 
    5493, 
    2512, 
    2923, 
    5984, 
    5483, 
    5676, 
    4010, 
    6232, 
    4239, 
    5536, 
    5715, 
    6513, 
    2804, 
    2512, 
    6391, 
    5829, 
    6249, 
    5651, 
    6028, 
    5602, 
    5765, 
    5546, 
    6208, 
    5724, 
    5765, 
    5602, 
    5779, 
    6338, 
    5904, 
    5617, 
    6028, 
    2923, 
    3265, 
    5904, 
    6459, 
    5765, 
    5493, 
    2923, 
    6028, 
    3265, 
    3573, 
    5602, 
    5984, 
    4450, 
    4239, 
    5483, 
    5984, 
    5573, 
    5676, 
    4450, 
    5984, 
    3897, 
    4450, 
    3629, 
    6232, 
    4010, 
    5940, 
    5536, 
    6232, 
    5940, 
    5573, 
    5984, 
    6232, 
    3897, 
    4239, 
    4450, 
    6014, 
    5806, 
    5090, 
    5715, 
    6014, 
    5219, 
    5715, 
    5536, 
    6014, 
    4955, 
    2523, 
    2932, 
    2552, 
    4955, 
    3629, 
    5264, 
    4539, 
    2523, 
    2552, 
    5264, 
    4955, 
    2552, 
    2956, 
    5264, 
    4701, 
    4872, 
    3580, 
    4734, 
    1504, 
    2771, 
    3458, 
    4734, 
    2771, 
    2528, 
    2418, 
    4734, 
    1005, 
    1782, 
    2609, 
    716, 
    4428, 
    6193, 
    4877, 
    851, 
    4533, 
    1175, 
    4877, 
    2200, 
    4331, 
    1664, 
    4877, 
    5427, 
    2008, 
    4494, 
    4331, 
    5130, 
    4986, 
    544, 
    2008, 
    5130, 
    1754, 
    1203, 
    1920, 
    4331, 
    4986, 
    1664, 
    851, 
    4877, 
    1664, 
    810, 
    544, 
    5130, 
    970, 
    1203, 
    1754, 
    543, 
    1179, 
    2008, 
    5105, 
    2549, 
    6305, 
    2060, 
    5105, 
    2819, 
    5072, 
    2549, 
    5105, 
    1705, 
    5072, 
    911, 
    3354, 
    4590, 
    5072, 
    2256, 
    3657, 
    1705, 
    4590, 
    2954, 
    2549, 
    2635, 
    4590, 
    3354, 
    2635, 
    1514, 
    4590, 
    851, 
    1664, 
    2426, 
    5795, 
    3490, 
    3775, 
    3349, 
    5795, 
    3015, 
    3349, 
    6194, 
    5795, 
    4598, 
    1671, 
    2229, 
    1911, 
    4598, 
    970, 
    1911, 
    1470, 
    4598, 
    861, 
    2035, 
    2465, 
    6170, 
    1048, 
    2138, 
    6170, 
    5531, 
    2659, 
    5001, 
    6170, 
    2138, 
    6517, 
    6068, 
    6451, 
    1546, 
    5001, 
    2138, 
    5944, 
    2608, 
    3331, 
    5656, 
    6451, 
    5809, 
    6106, 
    1371, 
    2033, 
    6068, 
    6106, 
    5944, 
    6068, 
    3825, 
    6106, 
    3945, 
    3046, 
    3675, 
    4203, 
    3949, 
    3678, 
    3380, 
    3046, 
    3411, 
    3973, 
    3678, 
    3708, 
    2465, 
    3973, 
    2882, 
    4203, 
    1373, 
    3949, 
    2465, 
    4203, 
    3973, 
    2465, 
    2035, 
    4203, 
    3376, 
    3675, 
    3380, 
    5531, 
    6422, 
    3043, 
    3675, 
    3046, 
    3380, 
    5870, 
    3675, 
    3376, 
    3043, 
    5870, 
    3376, 
    5656, 
    5554, 
    6369, 
    6231, 
    5554, 
    2605, 
    5122, 
    6231, 
    2605, 
    5814, 
    5949, 
    6369, 
    6422, 
    5656, 
    5870, 
    3043, 
    6422, 
    5870, 
    5531, 
    6170, 
    6517, 
    6517, 
    6170, 
    5001, 
    2994, 
    2605, 
    5554, 
    3945, 
    2664, 
    3046, 
    6369, 
    5554, 
    6231, 
    5122, 
    3806, 
    3527, 
    2664, 
    2706, 
    3082, 
    4981, 
    3215, 
    5972, 
    6382, 
    5949, 
    5814, 
    2664, 
    6382, 
    4370, 
    3945, 
    5949, 
    6382, 
    3527, 
    3215, 
    4981, 
    2366, 
    4082, 
    1845, 
    4391, 
    2706, 
    2664, 
    2166, 
    1095, 
    2706, 
    1809, 
    1048, 
    2659, 
    4680, 
    3678, 
    3949, 
    3043, 
    4680, 
    4501, 
    3043, 
    3376, 
    4680, 
    3547, 
    2343, 
    1373, 
    4904, 
    3547, 
    1373, 
    1889, 
    525, 
    4089, 
    3547, 
    4304, 
    2343, 
    4304, 
    4593, 
    1809, 
    4369, 
    4232, 
    4444, 
    2092, 
    4232, 
    1460, 
    3569, 
    3262, 
    4232, 
    2974, 
    3569, 
    956, 
    2974, 
    2581, 
    3569, 
    1188, 
    2092, 
    1460, 
    1188, 
    1095, 
    2220, 
    4300, 
    4000, 
    1412, 
    2366, 
    4300, 
    1412, 
    1140, 
    2191, 
    4300, 
    2220, 
    1660, 
    956, 
    1188, 
    2220, 
    2092, 
    1095, 
    2166, 
    2220, 
    1845, 
    1095, 
    1188, 
    2392, 
    1877, 
    1909, 
    1188, 
    2392, 
    1909, 
    5216, 
    5857, 
    3178, 
    2465, 
    2628, 
    861, 
    1909, 
    2366, 
    1845, 
    4449, 
    3775, 
    3490, 
    1920, 
    4449, 
    2954, 
    1203, 
    3775, 
    4449, 
    3172, 
    2819, 
    5105, 
    2954, 
    4449, 
    6305, 
    6180, 
    3230, 
    3540, 
    4082, 
    6180, 
    3540, 
    3652, 
    3349, 
    6180, 
    3490, 
    5795, 
    6194, 
    3015, 
    2882, 
    6190, 
    2882, 
    3015, 
    2628, 
    3817, 
    3082, 
    2706, 
    2366, 
    3924, 
    4082, 
    3230, 
    3411, 
    3540, 
    6190, 
    3230, 
    6180, 
    3015, 
    6190, 
    3349, 
    2882, 
    3230, 
    6190, 
    3708, 
    3380, 
    3411, 
    2882, 
    3708, 
    3230, 
    2882, 
    3973, 
    3708, 
    1412, 
    2060, 
    2819, 
    4203, 
    2035, 
    1373, 
    3411, 
    3230, 
    3708, 
    3082, 
    3411, 
    3046, 
    3082, 
    3540, 
    3411, 
    2664, 
    3082, 
    3046, 
    3817, 
    1095, 
    1845, 
    3082, 
    3817, 
    3540, 
    2706, 
    1095, 
    3817, 
    6194, 
    3349, 
    3652, 
    3172, 
    6194, 
    3652, 
    3172, 
    3490, 
    6194, 
    3852, 
    767, 
    1604, 
    1155, 
    3852, 
    831, 
    1155, 
    1986, 
    3852, 
    1664, 
    4986, 
    1754, 
    6020, 
    2635, 
    3657, 
    6494, 
    6020, 
    3657, 
    2256, 
    6494, 
    3657, 
    1242, 
    4526, 
    6494, 
    4526, 
    767, 
    6020, 
    1664, 
    1920, 
    2426, 
    2426, 
    2954, 
    4590, 
    851, 
    2426, 
    1514, 
    4590, 
    2549, 
    5072, 
    1920, 
    2954, 
    2426, 
    1920, 
    1203, 
    4449, 
    1473, 
    1038, 
    560, 
    2402, 
    1604, 
    1473, 
    1775, 
    2402, 
    1349, 
    1775, 
    831, 
    2402, 
    2325, 
    1038, 
    1473, 
    2102, 
    981, 
    1116, 
    1862, 
    2102, 
    1116, 
    4735, 
    1339, 
    2323, 
    1480, 
    4735, 
    2102, 
    1480, 
    2013, 
    4735, 
    2185, 
    1130, 
    2629, 
    5317, 
    2185, 
    2629, 
    818, 
    5317, 
    2013, 
    1613, 
    2185, 
    5317, 
    4888, 
    1253, 
    885, 
    1613, 
    4888, 
    2185, 
    5173, 
    1394, 
    1253, 
    1613, 
    5173, 
    4888, 
    1613, 
    779, 
    5173, 
    4600, 
    2388, 
    3388, 
    3685, 
    4600, 
    3388, 
    3499, 
    1870, 
    4600, 
    3782, 
    5429, 
    3499, 
    1130, 
    4006, 
    3016, 
    4079, 
    2424, 
    1512, 
    4835, 
    4079, 
    1512, 
    2117, 
    4835, 
    1512, 
    3502, 
    4659, 
    4835, 
    3815, 
    6270, 
    4079, 
    3937, 
    2278, 
    1275, 
    5003, 
    3815, 
    2461, 
    2879, 
    4954, 
    5003, 
    3854, 
    2525, 
    4800, 
    1732, 
    2278, 
    3276, 
    3024, 
    3731, 
    2195, 
    4437, 
    4079, 
    6270, 
    1918, 
    4437, 
    2933, 
    1918, 
    2424, 
    4437, 
    4294, 
    1732, 
    946, 
    2424, 
    4079, 
    4437, 
    4954, 
    5094, 
    3582, 
    3527, 
    3666, 
    3937, 
    3666, 
    3365, 
    3582, 
    3937, 
    3666, 
    3276, 
    2278, 
    3937, 
    3276, 
    1275, 
    3215, 
    3937, 
    3527, 
    3806, 
    3666, 
    5949, 
    3945, 
    3675, 
    5870, 
    5949, 
    3675, 
    5814, 
    4981, 
    6382, 
    6369, 
    6231, 
    5814, 
    5870, 
    6369, 
    5949, 
    5870, 
    5656, 
    6369, 
    5122, 
    4981, 
    5814, 
    3806, 
    5122, 
    2605, 
    4981, 
    4370, 
    6382, 
    5972, 
    4565, 
    4981, 
    1974, 
    5972, 
    3215, 
    1974, 
    747, 
    5972, 
    2664, 
    3945, 
    6382, 
    3806, 
    3365, 
    3666, 
    4981, 
    5122, 
    3527, 
    2605, 
    4068, 
    3806, 
    6270, 
    2525, 
    4437, 
    4800, 
    6270, 
    3815, 
    4800, 
    2525, 
    6270, 
    3365, 
    3854, 
    3582, 
    3033, 
    2525, 
    3854, 
    1034, 
    1799, 
    2278, 
    2227, 
    4177, 
    4495, 
    4219, 
    960, 
    876, 
    1918, 
    2638, 
    2424, 
    4887, 
    960, 
    4219, 
    4797, 
    4887, 
    4219, 
    3024, 
    2195, 
    4887, 
    4887, 
    2195, 
    960, 
    1918, 
    3024, 
    2638, 
    3731, 
    1625, 
    2195, 
    1201, 
    3731, 
    3024, 
    1201, 
    2227, 
    3731, 
    1625, 
    2316, 
    2195, 
    4306, 
    796, 
    1625, 
    2227, 
    4306, 
    3731, 
    2227, 
    1669, 
    4306, 
    1625, 
    3552, 
    2316, 
    6230, 
    6401, 
    4938, 
    5080, 
    467, 
    466, 
    3088, 
    5080, 
    1283, 
    3088, 
    1103, 
    5207, 
    3122, 
    3246, 
    1103, 
    1589, 
    473, 
    6120, 
    2085, 
    1450, 
    678, 
    2879, 
    2085, 
    946, 
    1732, 
    5094, 
    946, 
    4045, 
    3388, 
    1450, 
    2461, 
    4045, 
    2879, 
    2461, 
    3785, 
    4045, 
    5094, 
    3276, 
    3582, 
    2879, 
    5094, 
    4954, 
    1732, 
    3276, 
    5094, 
    4835, 
    2117, 
    3502, 
    1786, 
    3782, 
    3954, 
    6156, 
    4711, 
    1394, 
    5788, 
    4622, 
    4343, 
    5004, 
    4429, 
    4215, 
    5788, 
    4343, 
    4131, 
    5147, 
    4622, 
    4429, 
    5004, 
    5147, 
    4429, 
    1955, 
    716, 
    5147, 
    716, 
    1557, 
    4622, 
    6039, 
    5882, 
    2535, 
    6387, 
    6039, 
    2467, 
    3282, 
    6387, 
    2467, 
    3282, 
    5743, 
    6387, 
    6257, 
    2532, 
    2489, 
    6387, 
    6257, 
    6039, 
    5743, 
    2532, 
    6257, 
    4001, 
    1249, 
    1955, 
    716, 
    4622, 
    5147, 
    5165, 
    3089, 
    2262, 
    1249, 
    5165, 
    2262, 
    4227, 
    5028, 
    5165, 
    5004, 
    4227, 
    4001, 
    5147, 
    5004, 
    4001, 
    4215, 
    5495, 
    5004, 
    5028, 
    2733, 
    3415, 
    5495, 
    4441, 
    4227, 
    3988, 
    3724, 
    5538, 
    4804, 
    2733, 
    5538, 
    4958, 
    3103, 
    4804, 
    5098, 
    3722, 
    3432, 
    2736, 
    5098, 
    4958, 
    3818, 
    5478, 
    5098, 
    6108, 
    3818, 
    2736, 
    6328, 
    6258, 
    6377, 
    3106, 
    6328, 
    2736, 
    3106, 
    3435, 
    6339, 
    6393, 
    6260, 
    3541, 
    5621, 
    6393, 
    6108, 
    5621, 
    6441, 
    6393, 
    5478, 
    3987, 
    3722, 
    3541, 
    5478, 
    3818, 
    3541, 
    3232, 
    5585, 
    6464, 
    6203, 
    6293, 
    3987, 
    4213, 
    3556, 
    5596, 
    3256, 
    2748, 
    3711, 
    5596, 
    2748, 
    3976, 
    5366, 
    5596, 
    5366, 
    2501, 
    2524, 
    5596, 
    5366, 
    3256, 
    3976, 
    4205, 
    5366, 
    3103, 
    3976, 
    3711, 
    4205, 
    3722, 
    4095, 
    5366, 
    2524, 
    3256, 
    1249, 
    4001, 
    5165, 
    1712, 
    4536, 
    4880, 
    5816, 
    3853, 
    4119, 
    6075, 
    5816, 
    4119, 
    4711, 
    4544, 
    6466, 
    1394, 
    4711, 
    1253, 
    4544, 
    5739, 
    6466, 
    1394, 
    721, 
    6156, 
    6074, 
    4223, 
    3275, 
    4544, 
    6074, 
    5739, 
    2556, 
    4133, 
    6074, 
    6039, 
    2489, 
    5882, 
    6387, 
    5743, 
    6257, 
    1426, 
    1222, 
    2532, 
    6075, 
    1690, 
    885, 
    3838, 
    1456, 
    2389, 
    4536, 
    3838, 
    2389, 
    918, 
    2066, 
    3838, 
    2082, 
    710, 
    874, 
    1446, 
    2082, 
    874, 
    1305, 
    2296, 
    2082, 
    2082, 
    941, 
    710, 
    3480, 
    1456, 
    2089, 
    952, 
    4868, 
    4977, 
    4825, 
    4895, 
    4720, 
    5671, 
    2766, 
    5996, 
    4033, 
    5671, 
    3766, 
    4033, 
    1305, 
    6456, 
    2587, 
    4033, 
    3766, 
    1305, 
    5666, 
    6456, 
    2449, 
    2867, 
    5042, 
    3480, 
    4825, 
    1456, 
    4536, 
    1712, 
    918, 
    1874, 
    4536, 
    2389, 
    1874, 
    1135, 
    4880, 
    5304, 
    2449, 
    3129, 
    774, 
    5304, 
    3129, 
    1609, 
    1125, 
    6164, 
    1135, 
    3938, 
    4880, 
    1760, 
    975, 
    1726, 
    2283, 
    6267, 
    1739, 
    6267, 
    4868, 
    1739, 
    975, 
    6267, 
    4844, 
    4695, 
    4868, 
    6267, 
    1760, 
    4695, 
    975, 
    5422, 
    3766, 
    4977, 
    5739, 
    6074, 
    3581, 
    3853, 
    6466, 
    3581, 
    4544, 
    2556, 
    6074, 
    4223, 
    2501, 
    3275, 
    2066, 
    3564, 
    5414, 
    3564, 
    918, 
    3115, 
    3256, 
    3564, 
    2748, 
    2066, 
    918, 
    3564, 
    3115, 
    2748, 
    3564, 
    1712, 
    3115, 
    918, 
    3415, 
    2733, 
    3711, 
    3089, 
    3415, 
    3115, 
    5028, 
    4227, 
    4441, 
    2099, 
    465, 
    464, 
    1283, 
    1475, 
    2099, 
    1283, 
    466, 
    1475, 
    1726, 
    2274, 
    458, 
    6496, 
    2616, 
    6095, 
    5821, 
    6496, 
    6095, 
    1749, 
    1039, 
    6496, 
    5378, 
    4616, 
    6093, 
    1036, 
    1530, 
    2131, 
    5360, 
    2005, 
    800, 
    1205, 
    5360, 
    5155, 
    681, 
    2005, 
    5360, 
    2124, 
    681, 
    1205, 
    1241, 
    640, 
    366, 
    1241, 
    812, 
    367, 
    5308, 
    2058, 
    2880, 
    2058, 
    1352, 
    703, 
    5214, 
    2719, 
    2785, 
    5764, 
    6471, 
    2785, 
    2363, 
    1842, 
    5214, 
    908, 
    1352, 
    2058, 
    704, 
    5086, 
    3599, 
    4416, 
    1629, 
    890, 
    3007, 
    5822, 
    2495, 
    5378, 
    5155, 
    800, 
    4416, 
    5378, 
    1629, 
    4416, 
    4616, 
    5378, 
    5939, 
    5524, 
    3065, 
    3396, 
    5939, 
    3065, 
    3959, 
    5524, 
    5939, 
    3691, 
    3959, 
    5939, 
    2625, 
    704, 
    4191, 
    1842, 
    2719, 
    5214, 
    6521, 
    4071, 
    4290, 
    6283, 
    5568, 
    3368, 
    2585, 
    4071, 
    5568, 
    890, 
    1629, 
    4018, 
    3094, 
    2785, 
    2719, 
    3803, 
    2163, 
    3669, 
    4789, 
    2685, 
    3144, 
    5923, 
    4789, 
    3144, 
    2861, 
    2442, 
    4789, 
    2442, 
    2861, 
    2650, 
    5494, 
    3065, 
    2685, 
    2442, 
    5494, 
    4789, 
    2442, 
    4209, 
    5494, 
    4931, 
    1653, 
    1055, 
    2363, 
    4931, 
    1842, 
    4851, 
    834, 
    4931, 
    2363, 
    4851, 
    4931, 
    5821, 
    684, 
    965, 
    5638, 
    5369, 
    2753, 
    3120, 
    6113, 
    2753, 
    5454, 
    5344, 
    5638, 
    6171, 
    684, 
    5369, 
    5646, 
    1885, 
    4767, 
    3893, 
    3136, 
    3460, 
    3748, 
    5481, 
    3460, 
    2585, 
    6058, 
    3893, 
    5086, 
    371, 
    370, 
    2625, 
    2005, 
    1056, 
    812, 
    4407, 
    704, 
    5426, 
    2005, 
    2625, 
    3959, 
    5426, 
    2625, 
    3959, 
    3691, 
    5426, 
    372, 
    371, 
    1056, 
    1038, 
    562, 
    561, 
    560, 
    1038, 
    561, 
    4484, 
    2107, 
    1489, 
    6300, 
    4484, 
    3577, 
    562, 
    6300, 
    3577, 
    1038, 
    2325, 
    6300, 
    707, 
    4050, 
    4484, 
    930, 
    1718, 
    2112, 
    6402, 
    1018, 
    1359, 
    3343, 
    6402, 
    1359, 
    6242, 
    3469, 
    6402, 
    1344, 
    3105, 
    1029, 
    849, 
    2029, 
    3422, 
    2811, 
    1036, 
    841, 
    4413, 
    2811, 
    1519, 
    1802, 
    1036, 
    2811, 
    1359, 
    2722, 
    4413, 
    1931, 
    671, 
    1802, 
    2339, 
    1931, 
    1802, 
    4573, 
    701, 
    4167, 
    1931, 
    4573, 
    4167, 
    1217, 
    2236, 
    4775, 
    2131, 
    1205, 
    1656, 
    1036, 
    2131, 
    1656, 
    1530, 
    2124, 
    2131, 
    4080, 
    2727, 
    1530, 
    1931, 
    5865, 
    671, 
    1239, 
    377, 
    4080, 
    2124, 
    374, 
    681, 
    2727, 
    2124, 
    1530, 
    376, 
    375, 
    2124, 
    671, 
    1530, 
    1036, 
    2017, 
    1532, 
    826, 
    1650, 
    4703, 
    6094, 
    1344, 
    1532, 
    2017, 
    6242, 
    3343, 
    5960, 
    3147, 
    6242, 
    5960, 
    3469, 
    3756, 
    6286, 
    6289, 
    5643, 
    5798, 
    1984, 
    5964, 
    1294, 
    5485, 
    5678, 
    6528, 
    3915, 
    2530, 
    5156, 
    4163, 
    2937, 
    2530, 
    3585, 
    3278, 
    5523, 
    3083, 
    3857, 
    2707, 
    1029, 
    3756, 
    6011, 
    5576, 
    3756, 
    3469, 
    3278, 
    3998, 
    3734, 
    3278, 
    3585, 
    3998, 
    4886, 
    3469, 
    3147, 
    2789, 
    5037, 
    3147, 
    3734, 
    3998, 
    5576, 
    5615, 
    3734, 
    3446, 
    5907, 
    5615, 
    3446, 
    2937, 
    3734, 
    5615, 
    6011, 
    3585, 
    3857, 
    5576, 
    6011, 
    3756, 
    3998, 
    3585, 
    6011, 
    6095, 
    6390, 
    5821, 
    5425, 
    5454, 
    2620, 
    1885, 
    5344, 
    4377, 
    5344, 
    6171, 
    5638, 
    2909, 
    4416, 
    890, 
    1036, 
    1656, 
    841, 
    5378, 
    800, 
    1629, 
    4786, 
    6093, 
    4616, 
    1205, 
    681, 
    5360, 
    4191, 
    5524, 
    3959, 
    1056, 
    704, 
    2625, 
    5600, 
    3227, 
    2880, 
    2685, 
    5524, 
    6010, 
    6309, 
    4407, 
    5876, 
    6487, 
    6309, 
    5876, 
    5524, 
    4191, 
    6309, 
    363, 
    362, 
    1023, 
    5905, 
    6665, 
    1410, 
    1273, 
    5467, 
    3510, 
    4719, 
    5041, 
    4024, 
    6225, 
    969, 
    1403, 
    5601, 
    2563, 
    5590, 
    5601, 
    1298, 
    2563, 
    2194, 
    1526, 
    665, 
    2194, 
    1624, 
    1526, 
    2868, 
    3012, 
    1144, 
    2821, 
    5149, 
    3060, 
    4747, 
    2821, 
    1624, 
    3012, 
    4747, 
    2194, 
    3012, 
    3347, 
    4747, 
    1144, 
    3012, 
    2194, 
    4198, 
    5937, 
    3966, 
    3921, 
    3651, 
    6111, 
    1753, 
    4858, 
    969, 
    3776, 
    3651, 
    3921, 
    5590, 
    4716, 
    2680, 
    5601, 
    5590, 
    4858, 
    1753, 
    5601, 
    4858, 
    1082, 
    1298, 
    5601, 
    2563, 
    4716, 
    5590, 
    3492, 
    3347, 
    3776, 
    4747, 
    3347, 
    3492, 
    3012, 
    2450, 
    3347, 
    795, 
    2123, 
    1624, 
    3947, 
    944, 
    2583, 
    3242, 
    3947, 
    2178, 
    3242, 
    1730, 
    3947, 
    764, 
    4515, 
    5924, 
    4665, 
    3510, 
    3195, 
    4056, 
    4665, 
    4488, 
    2276, 
    3510, 
    4665, 
    3242, 
    2276, 
    1730, 
    944, 
    3947, 
    1730, 
    1600, 
    764, 
    5924, 
    3510, 
    2845, 
    3195, 
    4488, 
    4665, 
    3195, 
    1273, 
    1972, 
    5467, 
    4488, 
    1180, 
    1904, 
    1730, 
    4665, 
    4056, 
    3195, 
    1180, 
    4488, 
    3195, 
    2215, 
    1180, 
    1273, 
    3510, 
    2276, 
    2845, 
    1654, 
    3195, 
    1654, 
    5040, 
    4654, 
    5407, 
    5040, 
    837, 
    1180, 
    5515, 
    3204, 
    1654, 
    4654, 
    2215, 
    5515, 
    2854, 
    3204, 
    1082, 
    5515, 
    4654, 
    1082, 
    1753, 
    5515, 
    5515, 
    1753, 
    2854, 
    5358, 
    4909, 
    1903, 
    4044, 
    5358, 
    1177, 
    4044, 
    2693, 
    5358, 
    6126, 
    6395, 
    4314, 
    2832, 
    3964, 
    3698, 
    5537, 
    4314, 
    4098, 
    5716, 
    5537, 
    4462, 
    6557, 
    6301, 
    6463, 
    6301, 
    5898, 
    6215, 
    6371, 
    6463, 
    6215, 
    3620, 
    3889, 
    6301, 
    6312, 
    5533, 
    5756, 
    6420, 
    6215, 
    5878, 
    6126, 
    6550, 
    6013, 
    6463, 
    6301, 
    6215, 
    6550, 
    6463, 
    6371, 
    6372, 
    6550, 
    6371, 
    6126, 
    5537, 
    6550, 
    5716, 
    3313, 
    6557, 
    5527, 
    5533, 
    5883, 
    3889, 
    5898, 
    6301, 
    5709, 
    2798, 
    5457, 
    5537, 
    4098, 
    4462, 
    6013, 
    6550, 
    6372, 
    4196, 
    4270, 
    4314, 
    2832, 
    5464, 
    3964, 
    4270, 
    4098, 
    4314, 
    5390, 
    4270, 
    4196, 
    5464, 
    5390, 
    4196, 
    2634, 
    1928, 
    5390, 
    1212, 
    2234, 
    4270, 
    2234, 
    1680, 
    4098, 
    4126, 
    3990, 
    2926, 
    5951, 
    4126, 
    3862, 
    6423, 
    5951, 
    3862, 
    2538, 
    6423, 
    3862, 
    5532, 
    5033, 
    6423, 
    4881, 
    2602, 
    6502, 
    4538, 
    3330, 
    4339, 
    2225, 
    4655, 
    1197, 
    4655, 
    1867, 
    1124, 
    1197, 
    4655, 
    4578, 
    2225, 
    1369, 
    4690, 
    4690, 
    1867, 
    4655, 
    2411, 
    2519, 
    1445, 
    2519, 
    1867, 
    2384, 
    1445, 
    2519, 
    2384, 
    1489, 
    2107, 
    5320, 
    4110, 
    4324, 
    4697, 
    2107, 
    990, 
    4697, 
    3596, 
    1716, 
    925, 
    2934, 
    2526, 
    2554, 
    1541, 
    2934, 
    2554, 
    1541, 
    1336, 
    6274, 
    6138, 
    6274, 
    2636, 
    5108, 
    1541, 
    689, 
    6274, 
    1043, 
    2636, 
    2934, 
    6274, 
    6138, 
    1336, 
    1043, 
    6274, 
    1805, 
    4417, 
    2636, 
    6041, 
    1999, 
    4179, 
    2264, 
    6041, 
    4179, 
    4058, 
    1999, 
    6041, 
    2441, 
    830, 
    1744, 
    2286, 
    2441, 
    1744, 
    2286, 
    1652, 
    2441, 
    1980, 
    2212, 
    1289, 
    2910, 
    2496, 
    4034, 
    3526, 
    2860, 
    3210, 
    2445, 
    2496, 
    2846, 
    2962, 
    2410, 
    1488, 
    4466, 
    4258, 
    3005, 
    3646, 
    4648, 
    3341, 
    3252, 
    4258, 
    4466, 
    5151, 
    1595, 
    2175, 
    1901, 
    5151, 
    2410, 
    1901, 
    1595, 
    5151, 
    759, 
    1901, 
    1174, 
    5151, 
    2175, 
    5444, 
    3311, 
    4899, 
    5044, 
    5151, 
    5444, 
    2410, 
    759, 
    2674, 
    1595, 
    5444, 
    1488, 
    2410, 
    1108, 
    5444, 
    2175, 
    1108, 
    3851, 
    5444, 
    5242, 
    1174, 
    1901, 
    4277, 
    3791, 
    4051, 
    2212, 
    1174, 
    3162, 
    1289, 
    2212, 
    1652, 
    5242, 
    3162, 
    1174, 
    3741, 
    5242, 
    1901, 
    5127, 
    3162, 
    5242, 
    3303, 
    3452, 
    3741, 
    2764, 
    3005, 
    2618, 
    4023, 
    1832, 
    1077, 
    1893, 
    3758, 
    2837, 
    1158, 
    2203, 
    3758, 
    2154, 
    1077, 
    1637, 
    3187, 
    4364, 
    4561, 
    3187, 
    1077, 
    2154, 
    4067, 
    4286, 
    3383, 
    3051, 
    1259, 
    2806, 
    1333, 
    1962, 
    727, 
    2319, 
    1782, 
    1259, 
    1333, 
    2319, 
    1962, 
    3831, 
    3732, 
    3444, 
    1637, 
    3138, 
    3997, 
    1637, 
    2201, 
    3138, 
    1005, 
    2112, 
    1718, 
    3791, 
    830, 
    1652, 
    5971, 
    3051, 
    2806, 
    5382, 
    5971, 
    3481, 
    5382, 
    3383, 
    5971, 
    4286, 
    727, 
    1962, 
    978, 
    4067, 
    3383, 
    2100, 
    1477, 
    4869, 
    1962, 
    1259, 
    3051, 
    3791, 
    3511, 
    4491, 
    3880, 
    3519, 
    776, 
    4435, 
    3610, 
    3880, 
    1610, 
    4435, 
    3880, 
    2521, 
    3992, 
    4221, 
    5250, 
    5135, 
    3334, 
    3910, 
    5348, 
    3640, 
    3304, 
    2963, 
    5250, 
    2930, 
    3728, 
    3992, 
    5135, 
    4834, 
    2998, 
    3640, 
    5250, 
    3334, 
    2963, 
    2568, 
    5135, 
    3992, 
    3728, 
    3304, 
    3610, 
    4221, 
    3304, 
    2521, 
    2930, 
    3992, 
    4834, 
    2610, 
    2998, 
    3334, 
    5135, 
    2998, 
    2568, 
    4667, 
    4834, 
    3880, 
    3610, 
    3519, 
    1610, 
    3880, 
    776, 
    4474, 
    2183, 
    1127, 
    3610, 
    4435, 
    4221, 
    1610, 
    2183, 
    4435, 
    1307, 
    2805, 
    1990, 
    3285, 
    2266, 
    1718, 
    3481, 
    2806, 
    3285, 
    3767, 
    3481, 
    5459, 
    2298, 
    3767, 
    2805, 
    2298, 
    1762, 
    5382, 
    5382, 
    1762, 
    3383, 
    3051, 
    5971, 
    3383, 
    3767, 
    2298, 
    5382, 
    1259, 
    2266, 
    2806, 
    3468, 
    4458, 
    3146, 
    1962, 
    2319, 
    1259, 
    1566, 
    2009, 
    727, 
    6004, 
    3117, 
    2751, 
    6117, 
    6004, 
    2751, 
    3713, 
    4097, 
    6004, 
    5433, 
    3713, 
    2651, 
    5247, 
    5433, 
    2651, 
    5078, 
    2746, 
    5433, 
    4097, 
    3117, 
    6004, 
    3418, 
    4097, 
    3713, 
    3418, 
    3831, 
    4097, 
    3091, 
    3418, 
    2746, 
    3732, 
    3558, 
    3997, 
    3831, 
    3558, 
    3732, 
    3091, 
    2716, 
    3558, 
    2201, 
    1156, 
    3474, 
    3138, 
    2201, 
    3474, 
    4657, 
    4833, 
    5742, 
    2319, 
    4400, 
    1782, 
    4768, 
    3442, 
    3113, 
    4032, 
    4599, 
    3765, 
    4032, 
    4400, 
    4599, 
    1333, 
    3729, 
    2319, 
    1333, 
    2009, 
    3993, 
    5433, 
    2746, 
    3418, 
    3479, 
    4937, 
    3159, 
    4768, 
    3113, 
    4937, 
    3091, 
    3113, 
    2716, 
    4937, 
    5078, 
    6081, 
    4641, 
    3285, 
    1718, 
    4021, 
    4458, 
    3468, 
    4021, 
    2805, 
    4458, 
    1504, 
    2072, 
    930, 
    1433, 
    2378, 
    3843, 
    1504, 
    2418, 
    2072, 
    5539, 
    4610, 
    5498, 
    5834, 
    5539, 
    5498, 
    6414, 
    6280, 
    5498, 
    4412, 
    6414, 
    5498, 
    5610, 
    6280, 
    6414, 
    3316, 
    852, 
    5834, 
    5513, 
    5846, 
    5539, 
    1193, 
    4781, 
    5846, 
    1193, 
    2952, 
    4781, 
    5893, 
    4454, 
    1114, 
    852, 
    5893, 
    1114, 
    4730, 
    4553, 
    6373, 
    3073, 
    4730, 
    1599, 
    6373, 
    2780, 
    4454, 
    4730, 
    6373, 
    5893, 
    4553, 
    2780, 
    6373, 
    4357, 
    2780, 
    4553, 
    5440, 
    3208, 
    5279, 
    5047, 
    1868, 
    1127, 
    4454, 
    1859, 
    1114, 
    4015, 
    4245, 
    2780, 
    2595, 
    3843, 
    4922, 
    4922, 
    4245, 
    2595, 
    2378, 
    4922, 
    3843, 
    4454, 
    4245, 
    4922, 
    852, 
    1599, 
    5893, 
    2780, 
    4245, 
    4454, 
    3139, 
    5047, 
    4015, 
    2183, 
    2986, 
    3750, 
    2183, 
    1610, 
    3264, 
    3755, 
    1610, 
    776, 
    2378, 
    1193, 
    1859, 
    4454, 
    4922, 
    1859, 
    1433, 
    1912, 
    2378, 
    1599, 
    763, 
    3073, 
    5893, 
    1599, 
    4730, 
    2975, 
    2582, 
    5678, 
    5786, 
    2975, 
    5678, 
    763, 
    6220, 
    5485, 
    3316, 
    2975, 
    5786, 
    852, 
    3316, 
    6220, 
    4412, 
    4610, 
    3580, 
    4412, 
    3580, 
    3274, 
    5773, 
    6414, 
    4412, 
    5773, 
    5610, 
    6414, 
    3971, 
    6498, 
    4202, 
    6498, 
    4403, 
    6105, 
    4344, 
    2975, 
    6280, 
    5513, 
    852, 
    1114, 
    4610, 
    5539, 
    4781, 
    5539, 
    5834, 
    5513, 
    4731, 
    744, 
    1578, 
    5430, 
    5211, 
    1055, 
    2163, 
    5346, 
    4994, 
    2163, 
    1092, 
    5346, 
    4299, 
    3233, 
    4731, 
    5684, 
    5830, 
    1381, 
    3233, 
    744, 
    4731, 
    5081, 
    2470, 
    2887, 
    5629, 
    5856, 
    4993, 
    3748, 
    4127, 
    1749, 
    5856, 
    2539, 
    4993, 
    4127, 
    5856, 
    5629, 
    4336, 
    2539, 
    5856, 
    3460, 
    4336, 
    4127, 
    3460, 
    3136, 
    4336, 
    6058, 
    5374, 
    2776, 
    2978, 
    6058, 
    2585, 
    2978, 
    5374, 
    6058, 
    4987, 
    2275, 
    3591, 
    2886, 
    2859, 
    2438, 
    5629, 
    1294, 
    1039, 
    1749, 
    5629, 
    1039, 
    4127, 
    4336, 
    5856, 
    4535, 
    3136, 
    2776, 
    2539, 
    4535, 
    2944, 
    4336, 
    3136, 
    4535, 
    965, 
    3748, 
    1749, 
    4497, 
    6511, 
    1467, 
    4127, 
    3748, 
    3460, 
    965, 
    684, 
    6511, 
    4960, 
    3284, 
    3591, 
    1729, 
    4960, 
    3591, 
    4840, 
    5251, 
    4960, 
    2083, 
    4840, 
    943, 
    3208, 
    3520, 
    4840, 
    4336, 
    4535, 
    2539, 
    3591, 
    2275, 
    1729, 
    943, 
    4960, 
    1729, 
    6345, 
    2776, 
    4987, 
    3591, 
    6345, 
    4987, 
    3284, 
    4535, 
    6345, 
    4535, 
    3284, 
    2944, 
    4987, 
    1272, 
    2275, 
    3284, 
    6345, 
    3591, 
    2776, 
    3893, 
    6058, 
    2887, 
    2470, 
    4941, 
    1272, 
    2887, 
    2275, 
    1272, 
    1971, 
    3233, 
    3208, 
    2083, 
    1448, 
    5279, 
    3208, 
    1448, 
    2385, 
    5279, 
    1448, 
    4357, 
    5440, 
    5279, 
    3800, 
    3520, 
    2697, 
    3073, 
    3800, 
    2697, 
    5136, 
    2944, 
    5251, 
    4061, 
    5136, 
    3800, 
    2539, 
    2944, 
    5136, 
    5251, 
    3284, 
    4960, 
    4840, 
    2083, 
    3208, 
    689, 
    1940, 
    816, 
    2101, 
    979, 
    2669, 
    4243, 
    2101, 
    2669, 
    962, 
    4243, 
    2095, 
    962, 
    1478, 
    4243, 
    1478, 
    1400, 
    2101, 
    2051, 
    1400, 
    1478, 
    1693, 
    3980, 
    3320, 
    4725, 
    2175, 
    1595, 
    2674, 
    3953, 
    4725, 
    3311, 
    6071, 
    3627, 
    3902, 
    3634, 
    3953, 
    6071, 
    2982, 
    2589, 
    2971, 
    6071, 
    3311, 
    2971, 
    6182, 
    6071, 
    1833, 
    979, 
    2101, 
    5640, 
    3773, 
    4037, 
    4152, 
    5340, 
    2925, 
    4152, 
    3489, 
    5340, 
    1833, 
    2795, 
    1078, 
    4153, 
    2674, 
    759, 
    1289, 
    5185, 
    1980, 
    3902, 
    2674, 
    4153, 
    5185, 
    4653, 
    4470, 
    3634, 
    3684, 
    3953, 
    5160, 
    5379, 
    3902, 
    2514, 
    5640, 
    3326, 
    5456, 
    3327, 
    3634, 
    4037, 
    5456, 
    5379, 
    3773, 
    2795, 
    5456, 
    3327, 
    2774, 
    3684, 
    2990, 
    3327, 
    5456, 
    2990, 
    3055, 
    3327, 
    3834, 
    4862, 
    2196, 
    4783, 
    6057, 
    2824, 
    3239, 
    4613, 
    2898, 
    3239, 
    4414, 
    4613, 
    1883, 
    1146, 
    2482, 
    5435, 
    5287, 
    2395, 
    6333, 
    1308, 
    4244, 
    1883, 
    3251, 
    1146, 
    2299, 
    1308, 
    3251, 
    5287, 
    2299, 
    3251, 
    2395, 
    5287, 
    1883, 
    1763, 
    2299, 
    5287, 
    1763, 
    2155, 
    2299, 
    2155, 
    1567, 
    2299, 
    2989, 
    4470, 
    4653, 
    728, 
    1308, 
    1567, 
    1991, 
    777, 
    2788, 
    728, 
    1991, 
    1308, 
    728, 
    1963, 
    1991, 
    6000, 
    2228, 
    4085, 
    2219, 
    5143, 
    1186, 
    1202, 
    2228, 
    5143, 
    5060, 
    5228, 
    3603, 
    1894, 
    2405, 
    2288, 
    1159, 
    1894, 
    1292, 
    893, 
    2051, 
    2405, 
    1478, 
    962, 
    1747, 
    2405, 
    1478, 
    1747, 
    2356, 
    1833, 
    2101, 
    1400, 
    2356, 
    2101, 
    4550, 
    2577, 
    2971, 
    3055, 
    4550, 
    2774, 
    3055, 
    1400, 
    4550, 
    1833, 
    1078, 
    979, 
    5456, 
    4037, 
    3773, 
    3902, 
    5379, 
    3634, 
    4263, 
    4037, 
    5379, 
    5160, 
    4470, 
    4263, 
    4153, 
    5160, 
    3902, 
    5185, 
    1289, 
    4653, 
    4153, 
    5185, 
    5160, 
    4153, 
    1980, 
    5185, 
    3326, 
    5640, 
    4263, 
    1400, 
    2051, 
    4550, 
    3627, 
    2589, 
    3092, 
    1855, 
    3627, 
    3092, 
    3618, 
    3311, 
    3627, 
    4550, 
    2971, 
    5044, 
    6182, 
    3320, 
    2982, 
    2577, 
    6182, 
    2971, 
    2577, 
    3320, 
    6182, 
    5160, 
    4263, 
    5379, 
    2286, 
    4653, 
    1289, 
    2989, 
    3326, 
    4470, 
    3055, 
    2774, 
    3327, 
    2356, 
    3055, 
    2990, 
    2356, 
    1400, 
    3055, 
    759, 
    1980, 
    4153, 
    4244, 
    1991, 
    2788, 
    1627, 
    4244, 
    2788, 
    2196, 
    1146, 
    6333, 
    2856, 
    3834, 
    1627, 
    6333, 
    3251, 
    1308, 
    2196, 
    6333, 
    4244, 
    1146, 
    3251, 
    6333, 
    3518, 
    2436, 
    3206, 
    3551, 
    2342, 
    1372, 
    2034, 
    4414, 
    1372, 
    3239, 
    6269, 
    4316, 
    4862, 
    3834, 
    6269, 
    1808, 
    2342, 
    3551, 
    4244, 
    1308, 
    1991, 
    4862, 
    2898, 
    2482, 
    1146, 
    4862, 
    2482, 
    3834, 
    4100, 
    6269, 
    1627, 
    3834, 
    2196, 
    2856, 
    3206, 
    5496, 
    2315, 
    1808, 
    1047, 
    2196, 
    4862, 
    1146, 
    4316, 
    3551, 
    3239, 
    4414, 
    3551, 
    1372, 
    6057, 
    4613, 
    4414, 
    3176, 
    6057, 
    3939, 
    3176, 
    2824, 
    6057, 
    3239, 
    3551, 
    4414, 
    2990, 
    2795, 
    1833, 
    2356, 
    2990, 
    1833, 
    4725, 
    4899, 
    3618, 
    3327, 
    3684, 
    3634, 
    5044, 
    2971, 
    3311, 
    3684, 
    5044, 
    4899, 
    2774, 
    4550, 
    5044, 
    1308, 
    2299, 
    1567, 
    1763, 
    1078, 
    2155, 
    3251, 
    1883, 
    5287, 
    979, 
    1078, 
    1763, 
    4841, 
    1177, 
    1903, 
    1381, 
    6241, 
    1903, 
    4994, 
    1578, 
    2163, 
    6241, 
    4994, 
    4841, 
    4731, 
    1578, 
    4994, 
    5781, 
    6472, 
    4044, 
    1055, 
    5781, 
    4044, 
    1653, 
    4752, 
    6472, 
    5464, 
    2634, 
    5390, 
    3964, 
    5464, 
    4196, 
    3021, 
    2634, 
    5464, 
    5064, 
    4927, 
    3394, 
    3021, 
    5064, 
    4405, 
    5608, 
    4927, 
    5064, 
    3182, 
    5608, 
    5064, 
    3182, 
    3501, 
    5608, 
    3958, 
    2634, 
    3021, 
    664, 
    1928, 
    2634, 
    4994, 
    5346, 
    4841, 
    4462, 
    4098, 
    1680, 
    871, 
    4462, 
    1680, 
    3313, 
    5716, 
    4462, 
    4270, 
    5390, 
    1212, 
    1212, 
    5390, 
    1928, 
    5464, 
    2832, 
    3021, 
    5381, 
    5877, 
    6431, 
    3402, 
    3182, 
    3698, 
    5381, 
    6130, 
    5284, 
    3069, 
    3501, 
    3402, 
    5885, 
    2602, 
    4881, 
    5186, 
    5885, 
    5542, 
    5284, 
    6130, 
    5885, 
    4752, 
    1653, 
    834, 
    3394, 
    4927, 
    3063, 
    6141, 
    6472, 
    4752, 
    3069, 
    3784, 
    3501, 
    5781, 
    1055, 
    1653, 
    2693, 
    4044, 
    3784, 
    2693, 
    5680, 
    5358, 
    6472, 
    3784, 
    4044, 
    1653, 
    6472, 
    5781, 
    6141, 
    3784, 
    6472, 
    5186, 
    5542, 
    5054, 
    1177, 
    1055, 
    4044, 
    3063, 
    834, 
    703, 
    1352, 
    3920, 
    703, 
    3784, 
    3069, 
    2693, 
    6141, 
    3501, 
    3784, 
    4927, 
    6141, 
    4752, 
    4927, 
    5608, 
    6141, 
    3063, 
    4927, 
    4752, 
    3394, 
    3539, 
    5064, 
    3182, 
    3402, 
    3501, 
    6141, 
    5608, 
    3501, 
    3920, 
    3650, 
    3394, 
    703, 
    3920, 
    3063, 
    1352, 
    2745, 
    3920, 
    5064, 
    3021, 
    2832, 
    3539, 
    4405, 
    5064, 
    3539, 
    3229, 
    4405, 
    2832, 
    3698, 
    3182, 
    1928, 
    358, 
    1884, 
    2234, 
    4098, 
    4270, 
    664, 
    358, 
    1928, 
    4974, 
    5115, 
    2534, 
    5156, 
    5321, 
    3645, 
    5335, 
    5848, 
    6368, 
    5321, 
    6390, 
    3340, 
    6289, 
    1039, 
    5964, 
    6220, 
    3316, 
    5786, 
    5485, 
    6220, 
    5786, 
    1599, 
    852, 
    6220, 
    4202, 
    3274, 
    2932, 
    6105, 
    6099, 
    3587, 
    5773, 
    6105, 
    5610, 
    4403, 
    6099, 
    6105, 
    5513, 
    5834, 
    852, 
    4202, 
    5773, 
    4412, 
    6280, 
    3316, 
    5834, 
    3083, 
    673, 
    1532, 
    3857, 
    3083, 
    1532, 
    4028, 
    2779, 
    1219, 
    4271, 
    4254, 
    4047, 
    3083, 
    4271, 
    4047, 
    5523, 
    3278, 
    2937, 
    4479, 
    5523, 
    4376, 
    4479, 
    3585, 
    5523, 
    5226, 
    5376, 
    4645, 
    5271, 
    5174, 
    5097, 
    5371, 
    5271, 
    5226, 
    5323, 
    5371, 
    5226, 
    5628, 
    2679, 
    5328, 
    2558, 
    5628, 
    5371, 
    5790, 
    2894, 
    2478, 
    2558, 
    5790, 
    5628, 
    2558, 
    2757, 
    5981, 
    5328, 
    5229, 
    5174, 
    5628, 
    5328, 
    5271, 
    2679, 
    5312, 
    5328, 
    5452, 
    4254, 
    5376, 
    5097, 
    5452, 
    5376, 
    4957, 
    2779, 
    5452, 
    5328, 
    5312, 
    5229, 
    4803, 
    2779, 
    4957, 
    4047, 
    4254, 
    4028, 
    6514, 
    4163, 
    3915, 
    6514, 
    5522, 
    4163, 
    6326, 
    6514, 
    3915, 
    6326, 
    5579, 
    6514, 
    4974, 
    4821, 
    5522, 
    6210, 
    4821, 
    4974, 
    2534, 
    6210, 
    4974, 
    2757, 
    5323, 
    6210, 
    4645, 
    5852, 
    6091, 
    4742, 
    4479, 
    5852, 
    4254, 
    4742, 
    4464, 
    4271, 
    4479, 
    4742, 
    4479, 
    2707, 
    3585, 
    5852, 
    4479, 
    4376, 
    6091, 
    5852, 
    4376, 
    4645, 
    4464, 
    5852, 
    4271, 
    2707, 
    4479, 
    5523, 
    4163, 
    4376, 
    4254, 
    5452, 
    4028, 
    3233, 
    5081, 
    1272, 
    3820, 
    2470, 
    3543, 
    1679, 
    2886, 
    868, 
    1679, 
    2859, 
    2886, 
    4941, 
    1729, 
    2275, 
    6103, 
    4941, 
    2470, 
    2438, 
    6103, 
    2470, 
    2438, 
    5075, 
    6103, 
    2438, 
    5990, 
    5075, 
    5251, 
    4840, 
    3520, 
    3800, 
    5251, 
    3520, 
    2944, 
    3284, 
    5251, 
    4960, 
    943, 
    4840, 
    6511, 
    4497, 
    5481, 
    3748, 
    6511, 
    5481, 
    684, 
    1467, 
    6511, 
    5485, 
    1984, 
    763, 
    5678, 
    5485, 
    5786, 
    6368, 
    5678, 
    2582, 
    5643, 
    6528, 
    5678, 
    3587, 
    5335, 
    6368, 
    6289, 
    2616, 
    1039, 
    6528, 
    6289, 
    5964, 
    5485, 
    6528, 
    5964, 
    5643, 
    6289, 
    6528, 
    5798, 
    2616, 
    6289, 
    5964, 
    1984, 
    5485, 
    1749, 
    4127, 
    5629, 
    2616, 
    6496, 
    1039, 
    3136, 
    3893, 
    2776, 
    6345, 
    4535, 
    2776, 
    5646, 
    1467, 
    1226, 
    1885, 
    5646, 
    1226, 
    6511, 
    3748, 
    965, 
    4290, 
    5481, 
    4497, 
    4290, 
    6026, 
    5481, 
    5953, 
    4290, 
    4497, 
    3036, 
    6521, 
    2650, 
    6521, 
    5568, 
    4071, 
    2650, 
    6521, 
    5953, 
    3036, 
    5568, 
    6521, 
    6026, 
    3893, 
    5481, 
    4071, 
    6026, 
    4290, 
    4071, 
    2585, 
    6026, 
    2558, 
    5323, 
    2757, 
    2530, 
    3915, 
    4163, 
    5115, 
    2940, 
    2534, 
    5522, 
    5579, 
    4974, 
    5798, 
    6437, 
    3003, 
    5238, 
    5753, 
    5335, 
    6326, 
    3645, 
    5588, 
    5753, 
    6326, 
    5588, 
    5579, 
    5522, 
    6514, 
    5156, 
    3645, 
    3915, 
    5907, 
    5156, 
    2530, 
    5615, 
    5907, 
    2530, 
    6306, 
    5480, 
    5321, 
    3120, 
    6306, 
    5907, 
    3120, 
    2753, 
    6306, 
    6306, 
    2753, 
    6298, 
    5238, 
    3281, 
    2940, 
    5579, 
    5238, 
    5115, 
    4974, 
    5579, 
    5115, 
    3645, 
    3340, 
    5588, 
    5798, 
    3003, 
    2616, 
    5848, 
    6437, 
    5643, 
    6437, 
    3340, 
    3003, 
    5643, 
    6437, 
    5798, 
    5588, 
    3340, 
    6437, 
    5238, 
    2940, 
    5115, 
    5335, 
    3281, 
    5238, 
    6280, 
    5834, 
    5498, 
    4344, 
    6280, 
    5610, 
    2975, 
    3316, 
    6280, 
    4189, 
    3407, 
    3956, 
    4403, 
    3705, 
    4189, 
    6498, 
    6105, 
    5773, 
    4202, 
    6498, 
    5773, 
    3971, 
    4403, 
    6498, 
    2582, 
    4344, 
    3587, 
    2582, 
    2975, 
    4344, 
    2932, 
    2523, 
    3971, 
    2523, 
    4955, 
    5264, 
    3956, 
    3407, 
    3078, 
    5774, 
    3956, 
    3688, 
    5981, 
    5774, 
    3688, 
    3299, 
    3605, 
    5774, 
    4189, 
    3705, 
    3407, 
    5774, 
    5969, 
    3956, 
    6099, 
    3281, 
    3587, 
    3956, 
    5969, 
    4189, 
    3605, 
    3281, 
    6099, 
    6105, 
    3587, 
    4344, 
    4189, 
    6099, 
    4403, 
    5969, 
    3605, 
    6099, 
    4708, 
    5693, 
    4438, 
    3705, 
    4539, 
    3407, 
    3705, 
    2523, 
    4539, 
    5790, 
    3688, 
    2894, 
    3688, 
    3956, 
    3078, 
    2940, 
    3605, 
    3299, 
    5610, 
    6105, 
    4344, 
    3705, 
    4403, 
    3971, 
    4189, 
    5969, 
    6099, 
    5693, 
    4539, 
    5264, 
    2591, 
    5693, 
    2956, 
    4708, 
    4539, 
    5693, 
    2724, 
    5887, 
    4438, 
    3078, 
    3407, 
    4708, 
    4993, 
    4061, 
    1984, 
    5629, 
    4993, 
    1294, 
    2539, 
    5136, 
    4993, 
    3800, 
    5136, 
    5251, 
    992, 
    1773, 
    1679, 
    3177, 
    5315, 
    2825, 
    3257, 
    5389, 
    5463, 
    794, 
    1623, 
    1523, 
    2001, 
    794, 
    2430, 
    4102, 
    4318, 
    3421, 
    5796, 
    2475, 
    2926, 
    2497, 
    3969, 
    2911, 
    4356, 
    3224, 
    3536, 
    2891, 
    5258, 
    5353, 
    4145, 
    3224, 
    4356, 
    4969, 
    2875, 
    2458, 
    2756, 
    2737, 
    5327, 
    1320, 
    3056, 
    2001, 
    3095, 
    2309, 
    1773, 
    6311, 
    3421, 
    2538, 
    6311, 
    3267, 
    3421, 
    3862, 
    6311, 
    2538, 
    3862, 
    3267, 
    6311, 
    5532, 
    6423, 
    2538, 
    6502, 
    2992, 
    4538, 
    2926, 
    2475, 
    3836, 
    4318, 
    2309, 
    3095, 
    4902, 
    4075, 
    794, 
    2676, 
    4902, 
    3056, 
    4729, 
    4075, 
    4902, 
    1320, 
    2309, 
    4318, 
    2193, 
    1623, 
    2557, 
    3149, 
    2762, 
    2791, 
    2121, 
    2193, 
    1143, 
    1623, 
    794, 
    4075, 
    2121, 
    1623, 
    2193, 
    2379, 
    4453, 
    4889, 
    4639, 
    4216, 
    3989, 
    3317, 
    4889, 
    4712, 
    2379, 
    1434, 
    4453, 
    3056, 
    4902, 
    2001, 
    1860, 
    1115, 
    2583, 
    2976, 
    3389, 
    1115, 
    5924, 
    2276, 
    3242, 
    1600, 
    5924, 
    3242, 
    4515, 
    2276, 
    5924, 
    2976, 
    1115, 
    1860, 
    4889, 
    2976, 
    1860, 
    2379, 
    4889, 
    1860, 
    4453, 
    4712, 
    4889, 
    4889, 
    3317, 
    2976, 
    4639, 
    4712, 
    4453, 
    4639, 
    4545, 
    4712, 
    2875, 
    4145, 
    2458, 
    3702, 
    3404, 
    3686, 
    4855, 
    3702, 
    3686, 
    3317, 
    4855, 
    3686, 
    3623, 
    3891, 
    5758, 
    4790, 
    2739, 
    4946, 
    2497, 
    4790, 
    3702, 
    2497, 
    5594, 
    4790, 
    3404, 
    3075, 
    3389, 
    2976, 
    3686, 
    3389, 
    3702, 
    4790, 
    5987, 
    3075, 
    1600, 
    2178, 
    3389, 
    3075, 
    2178, 
    3317, 
    3686, 
    2976, 
    5758, 
    4855, 
    3623, 
    4145, 
    6332, 
    3891, 
    3969, 
    4855, 
    5758, 
    3389, 
    3686, 
    3404, 
    3317, 
    3623, 
    4855, 
    5092, 
    2739, 
    4630, 
    4951, 
    5092, 
    4442, 
    4946, 
    2739, 
    5092, 
    3404, 
    4946, 
    3075, 
    5987, 
    4790, 
    4946, 
    3404, 
    5987, 
    4946, 
    3404, 
    3702, 
    5987, 
    3242, 
    2178, 
    1600, 
    3947, 
    2583, 
    1115, 
    5330, 
    2386, 
    1449, 
    1774, 
    4373, 
    996, 
    3911, 
    1869, 
    4373, 
    2584, 
    1449, 
    2386, 
    3589, 
    2584, 
    2386, 
    2379, 
    5117, 
    2584, 
    4333, 
    4124, 
    2791, 
    1860, 
    5117, 
    2379, 
    2084, 
    5175, 
    1449, 
    5117, 
    2583, 
    2084, 
    2584, 
    5117, 
    1449, 
    1860, 
    2583, 
    5117, 
    944, 
    4393, 
    2084, 
    4056, 
    4488, 
    1904, 
    2412, 
    5373, 
    1904, 
    1730, 
    2276, 
    4665, 
    4515, 
    1273, 
    2276, 
    1985, 
    4515, 
    764, 
    1985, 
    4443, 
    4515, 
    2845, 
    837, 
    1654, 
    2215, 
    3195, 
    1654, 
    4976, 
    745, 
    4182, 
    3946, 
    4976, 
    4182, 
    4823, 
    2845, 
    5467, 
    2596, 
    1128, 
    4749, 
    2379, 
    2584, 
    1434, 
    3911, 
    4373, 
    1774, 
    3589, 
    2386, 
    1869, 
    2596, 
    3589, 
    1869, 
    1434, 
    2584, 
    3589, 
    5330, 
    2108, 
    996, 
    2386, 
    5330, 
    4373, 
    1449, 
    5175, 
    5330, 
    5175, 
    5895, 
    5330, 
    5175, 
    5373, 
    1494, 
    1730, 
    4393, 
    944, 
    4056, 
    1904, 
    5373, 
    1730, 
    4056, 
    4393, 
    2854, 
    1753, 
    969, 
    6225, 
    2854, 
    969, 
    4024, 
    6225, 
    1403, 
    4024, 
    3204, 
    6225, 
    1180, 
    3204, 
    1904, 
    1180, 
    4654, 
    5515, 
    1180, 
    2215, 
    4654, 
    4719, 
    4024, 
    1403, 
    2807, 
    4719, 
    2053, 
    5041, 
    1494, 
    2412, 
    2807, 
    5041, 
    4719, 
    2807, 
    5288, 
    5041, 
    5373, 
    4393, 
    4056, 
    1494, 
    5373, 
    2412, 
    5175, 
    4393, 
    5373, 
    5895, 
    5175, 
    1494, 
    2108, 
    5895, 
    1494, 
    2108, 
    5330, 
    5895, 
    2084, 
    4393, 
    5175, 
    1904, 
    3204, 
    4024, 
    2248, 
    1152, 
    1234, 
    4282, 
    3301, 
    3607, 
    1697, 
    1888, 
    2248, 
    3266, 
    728, 
    1567, 
    4439, 
    3266, 
    2925, 
    4225, 
    728, 
    3266, 
    3890, 
    2973, 
    3314, 
    2540, 
    3890, 
    3621, 
    4230, 
    3633, 
    3901, 
    5831, 
    4230, 
    4005, 
    6479, 
    5831, 
    4005, 
    3740, 
    6479, 
    4005, 
    5869, 
    4551, 
    6479, 
    4144, 
    4230, 
    5831, 
    2540, 
    3633, 
    4230, 
    1260, 
    777, 
    1963, 
    4807, 
    1611, 
    2267, 
    4749, 
    2184, 
    4807, 
    3563, 
    1324, 
    2004, 
    1128, 
    3563, 
    2184, 
    6268, 
    3911, 
    2312, 
    1128, 
    6268, 
    3563, 
    1128, 
    3911, 
    6268, 
    777, 
    1991, 
    1963, 
    1127, 
    3750, 
    5047, 
    4015, 
    2780, 
    3139, 
    2986, 
    4015, 
    3750, 
    2595, 
    4245, 
    4015, 
    4730, 
    3073, 
    2697, 
    3578, 
    3112, 
    3441, 
    3496, 
    3578, 
    3272, 
    3496, 
    2121, 
    3578, 
    2385, 
    3840, 
    5315, 
    3840, 
    1448, 
    2977, 
    4015, 
    2986, 
    2595, 
    5047, 
    3750, 
    4015, 
    3463, 
    5047, 
    3139, 
    3463, 
    1868, 
    5047, 
    1127, 
    2183, 
    3750, 
    3892, 
    3624, 
    3140, 
    1926, 
    3892, 
    3140, 
    2430, 
    3566, 
    3892, 
    3566, 
    3257, 
    3892, 
    3624, 
    2781, 
    3140, 
    5853, 
    3624, 
    3257, 
    2915, 
    5853, 
    3257, 
    2915, 
    2503, 
    5897, 
    3318, 
    2781, 
    3624, 
    2915, 
    5897, 
    5853, 
    2977, 
    5178, 
    5453, 
    5897, 
    2977, 
    3318, 
    5315, 
    3840, 
    2503, 
    2825, 
    5315, 
    2503, 
    3177, 
    1868, 
    5315, 
    2385, 
    1448, 
    3840, 
    1448, 
    2083, 
    2977, 
    5990, 
    2859, 
    4765, 
    2430, 
    794, 
    1523, 
    2430, 
    1926, 
    2001, 
    3566, 
    2430, 
    1523, 
    3496, 
    3566, 
    1523, 
    3257, 
    3624, 
    3892, 
    3624, 
    5853, 
    3318, 
    2121, 
    3496, 
    1523, 
    3496, 
    3272, 
    5389, 
    3566, 
    3496, 
    5389, 
    2121, 
    1022, 
    3578, 
    5897, 
    3840, 
    2977, 
    5853, 
    5897, 
    3318, 
    2503, 
    3840, 
    5897, 
    5203, 
    4941, 
    6103, 
    943, 
    5203, 
    5178, 
    943, 
    1729, 
    5203, 
    1209, 
    1320, 
    1926, 
    3264, 
    2986, 
    2183, 
    3755, 
    3264, 
    1610, 
    1990, 
    3755, 
    776, 
    3468, 
    5901, 
    3755, 
    5901, 
    3571, 
    3264, 
    3755, 
    5901, 
    3264, 
    3468, 
    3571, 
    5901, 
    3843, 
    2595, 
    3571, 
    3468, 
    4020, 
    3571, 
    2378, 
    1859, 
    4922, 
    4474, 
    2521, 
    4221, 
    2183, 
    4474, 
    4435, 
    3177, 
    2521, 
    4474, 
    3177, 
    2825, 
    2521, 
    1868, 
    3177, 
    1127, 
    1868, 
    2385, 
    5315, 
    2503, 
    2915, 
    5463, 
    1127, 
    3177, 
    4474, 
    4020, 
    2072, 
    1433, 
    2986, 
    3264, 
    3571, 
    4021, 
    3755, 
    1990, 
    5459, 
    4458, 
    2805, 
    3767, 
    5459, 
    2805, 
    3285, 
    4641, 
    5459, 
    3468, 
    3755, 
    4021, 
    4020, 
    3468, 
    3146, 
    4020, 
    3843, 
    3571, 
    2072, 
    4020, 
    3146, 
    1433, 
    3843, 
    4020, 
    2595, 
    2986, 
    3571, 
    4021, 
    1990, 
    2805, 
    763, 
    4061, 
    3073, 
    5453, 
    2781, 
    3318, 
    2977, 
    5453, 
    3318, 
    5075, 
    5990, 
    5453, 
    5178, 
    5075, 
    5453, 
    2083, 
    5178, 
    2977, 
    2083, 
    943, 
    5178, 
    5203, 
    6103, 
    5075, 
    4061, 
    763, 
    1984, 
    4061, 
    3800, 
    3073, 
    1294, 
    4993, 
    1984, 
    4993, 
    5136, 
    4061, 
    5893, 
    6373, 
    4454, 
    2697, 
    4553, 
    4730, 
    2697, 
    5440, 
    4553, 
    5279, 
    3463, 
    4357, 
    3463, 
    2385, 
    1868, 
    4357, 
    3463, 
    3139, 
    2780, 
    4357, 
    3139, 
    5440, 
    3520, 
    3208, 
    4553, 
    5440, 
    4357, 
    2697, 
    3520, 
    5440, 
    5279, 
    2385, 
    3463, 
    1799, 
    757, 
    2337, 
    5751, 
    5547, 
    6427, 
    3232, 
    5751, 
    2535, 
    6393, 
    3541, 
    3818, 
    5751, 
    6260, 
    6160, 
    3232, 
    3541, 
    6260, 
    4924, 
    4674, 
    4847, 
    5872, 
    4750, 
    5778, 
    4158, 
    6486, 
    3909, 
    6486, 
    4750, 
    5872, 
    4575, 
    4498, 
    4750, 
    6238, 
    3282, 
    2467, 
    3333, 
    5487, 
    3639, 
    3333, 
    2997, 
    5487, 
    5824, 
    3282, 
    6238, 
    3860, 
    3588, 
    5487, 
    1106, 
    3860, 
    2997, 
    1106, 
    1536, 
    3860, 
    5528, 
    1536, 
    678, 
    6421, 
    5528, 
    678, 
    5743, 
    6421, 
    1426, 
    5743, 
    5528, 
    6421, 
    2489, 
    6039, 
    6257, 
    3282, 
    3588, 
    5743, 
    3993, 
    3248, 
    2716, 
    3729, 
    3993, 
    3442, 
    3729, 
    1333, 
    3993, 
    2266, 
    1259, 
    1782, 
    1718, 
    2266, 
    1005, 
    3767, 
    5382, 
    3481, 
    4641, 
    4458, 
    5459, 
    2072, 
    4641, 
    930, 
    3146, 
    4458, 
    4641, 
    2072, 
    3146, 
    4641, 
    1307, 
    2298, 
    2805, 
    3383, 
    1762, 
    978, 
    2100, 
    4067, 
    978, 
    5971, 
    2806, 
    3481, 
    3285, 
    5459, 
    3481, 
    2266, 
    3285, 
    2806, 
    1718, 
    930, 
    4641, 
    5832, 
    3523, 
    3802, 
    2568, 
    4834, 
    5135, 
    4283, 
    3511, 
    2445, 
    5497, 
    4283, 
    4063, 
    6044, 
    5497, 
    4063, 
    2610, 
    4283, 
    5497, 
    4491, 
    2018, 
    830, 
    2610, 
    4372, 
    4283, 
    2610, 
    4658, 
    4372, 
    6227, 
    2997, 
    5517, 
    1593, 
    6227, 
    5517, 
    1034, 
    4294, 
    6227, 
    5824, 
    5487, 
    3588, 
    3282, 
    5824, 
    3588, 
    5544, 
    5722, 
    5824, 
    6238, 
    5544, 
    5824, 
    5751, 
    6427, 
    2467, 
    6427, 
    6019, 
    5544, 
    2467, 
    6427, 
    6238, 
    5547, 
    6019, 
    6427, 
    2535, 
    5751, 
    2467, 
    6042, 
    5689, 
    5696, 
    5722, 
    5862, 
    3639, 
    6019, 
    5722, 
    5544, 
    6238, 
    6427, 
    5544, 
    5696, 
    5511, 
    6019, 
    5862, 
    3909, 
    3639, 
    6137, 
    6001, 
    5890, 
    6019, 
    6137, 
    5722, 
    6019, 
    5511, 
    6137, 
    5890, 
    4158, 
    3909, 
    5722, 
    6137, 
    5862, 
    6115, 
    5620, 
    6086, 
    4158, 
    6115, 
    4371, 
    6001, 
    5620, 
    6115, 
    5862, 
    6137, 
    5890, 
    5511, 
    5620, 
    6001, 
    4847, 
    2951, 
    1979, 
    4847, 
    4674, 
    2951, 
    1593, 
    5061, 
    757, 
    5061, 
    5517, 
    5778, 
    4847, 
    5061, 
    4924, 
    1593, 
    1034, 
    6227, 
    4498, 
    3291, 
    4674, 
    2997, 
    3860, 
    5487, 
    5778, 
    3639, 
    5872, 
    5528, 
    3860, 
    1536, 
    2716, 
    3113, 
    3442, 
    2266, 
    1782, 
    1005, 
    3248, 
    3993, 
    2009, 
    3993, 
    2716, 
    3442, 
    811, 
    3248, 
    2009, 
    3997, 
    3138, 
    3732, 
    811, 
    3997, 
    3248, 
    811, 
    1637, 
    3997, 
    4723, 
    2956, 
    2552, 
    3479, 
    4768, 
    4937, 
    5247, 
    2651, 
    5742, 
    2804, 
    5247, 
    4833, 
    5078, 
    5433, 
    5247, 
    6081, 
    5078, 
    5247, 
    3159, 
    6081, 
    2804, 
    3159, 
    4937, 
    6081, 
    4937, 
    2746, 
    5078, 
    3732, 
    3138, 
    2778, 
    3444, 
    3732, 
    2778, 
    3558, 
    3248, 
    3997, 
    4833, 
    4657, 
    2923, 
    6081, 
    5247, 
    2804, 
    5742, 
    3037, 
    6344, 
    5247, 
    5742, 
    4833, 
    2651, 
    3037, 
    5742, 
    5056, 
    1065, 
    2936, 
    4914, 
    2352, 
    1822, 
    986, 
    4914, 
    1767, 
    986, 
    2906, 
    4914, 
    2771, 
    1504, 
    2112, 
    5022, 
    3274, 
    4872, 
    3705, 
    3971, 
    2523, 
    4557, 
    3747, 
    4360, 
    4529, 
    2952, 
    2528, 
    4734, 
    3458, 
    4557, 
    1114, 
    1859, 
    5846, 
    4557, 
    3458, 
    3747, 
    4529, 
    4557, 
    4360, 
    2528, 
    4734, 
    4557, 
    3274, 
    4202, 
    4412, 
    3971, 
    4202, 
    2932, 
    5846, 
    5513, 
    1114, 
    1193, 
    5846, 
    1859, 
    4781, 
    5539, 
    5846, 
    3580, 
    4610, 
    3292, 
    4412, 
    5498, 
    4610, 
    1193, 
    1912, 
    2952, 
    2418, 
    1504, 
    4734, 
    5056, 
    4914, 
    1822, 
    4222, 
    4211, 
    2747, 
    5110, 
    4970, 
    4890, 
    5174, 
    5229, 
    5038, 
    5084, 
    4970, 
    5110, 
    3994, 
    5084, 
    4222, 
    4944, 
    4970, 
    5084, 
    3730, 
    4944, 
    3994, 
    5110, 
    4890, 
    5038, 
    2044, 
    4970, 
    4944, 
    2044, 
    880, 
    4970, 
    4436, 
    3982, 
    4211, 
    5229, 
    5110, 
    5038, 
    5271, 
    5328, 
    5174, 
    5210, 
    5110, 
    5229, 
    4222, 
    5210, 
    4436, 
    5084, 
    5110, 
    5210, 
    6321, 
    2478, 
    4799, 
    4626, 
    3982, 
    4436, 
    5210, 
    5312, 
    4436, 
    6174, 
    3424, 
    4132, 
    3982, 
    6174, 
    3445, 
    4799, 
    3424, 
    6174, 
    6321, 
    4799, 
    4626, 
    2478, 
    2894, 
    4953, 
    3118, 
    2752, 
    4211, 
    2955, 
    2969, 
    3309, 
    2574, 
    4467, 
    4885, 
    3292, 
    4610, 
    4781, 
    5035, 
    2869, 
    2451, 
    4787, 
    4883, 
    4618, 
    4707, 
    2869, 
    4883, 
    3809, 
    3179, 
    3498, 
    2931, 
    3809, 
    3532, 
    2931, 
    3273, 
    3809, 
    6239, 
    3845, 
    3573, 
    5564, 
    6239, 
    3573, 
    4268, 
    4042, 
    6239, 
    3219, 
    4042, 
    2869, 
    3780, 
    5906, 
    6135, 
    3532, 
    3780, 
    3219, 
    3498, 
    5754, 
    5906, 
    3532, 
    3498, 
    3780, 
    4707, 
    3532, 
    3219, 
    2522, 
    2931, 
    3532, 
    5547, 
    5696, 
    6019, 
    5862, 
    5890, 
    3909, 
    3639, 
    5487, 
    5722, 
    6562, 
    6349, 
    6519, 
    5511, 
    5689, 
    5835, 
    6556, 
    5784, 
    5621, 
    6378, 
    6376, 
    6543, 
    5621, 
    6442, 
    6556, 
    6377, 
    6376, 
    6378, 
    6442, 
    6377, 
    6378, 
    6108, 
    6442, 
    5621, 
    6108, 
    6328, 
    6442, 
    6258, 
    6158, 
    6377, 
    6481, 
    6475, 
    5810, 
    6543, 
    6481, 
    6375, 
    6364, 
    6475, 
    6481, 
    5499, 
    5784, 
    5945, 
    5499, 
    6042, 
    6160, 
    5754, 
    6272, 
    4522, 
    6272, 
    2828, 
    5997, 
    5997, 
    2828, 
    4575, 
    4371, 
    5997, 
    4158, 
    4371, 
    6272, 
    5997, 
    6480, 
    5620, 
    5835, 
    4522, 
    6086, 
    6329, 
    4522, 
    4371, 
    6086, 
    6115, 
    4158, 
    5890, 
    6134, 
    5999, 
    6237, 
    3724, 
    6134, 
    3435, 
    6237, 
    5644, 
    6200, 
    6260, 
    5751, 
    3232, 
    6441, 
    6160, 
    6260, 
    5784, 
    6441, 
    5621, 
    5784, 
    5499, 
    6441, 
    6042, 
    5547, 
    6160, 
    6276, 
    6258, 
    6339, 
    6237, 
    6276, 
    6134, 
    6158, 
    6258, 
    6276, 
    6366, 
    6490, 
    6040, 
    6378, 
    6543, 
    6375, 
    6481, 
    5810, 
    5945, 
    6353, 
    6475, 
    6364, 
    6353, 
    6519, 
    6475, 
    6339, 
    6328, 
    3106, 
    6134, 
    6339, 
    3435, 
    6258, 
    6328, 
    6339, 
    6556, 
    6378, 
    6375, 
    5784, 
    6556, 
    6375, 
    6442, 
    6378, 
    6556, 
    6490, 
    6376, 
    6158, 
    6040, 
    6490, 
    6158, 
    6366, 
    6540, 
    6560, 
    6540, 
    6461, 
    6365, 
    6108, 
    2736, 
    6328, 
    6135, 
    4112, 
    3845, 
    6239, 
    6135, 
    3845, 
    4042, 
    3780, 
    6135, 
    3818, 
    6108, 
    6393, 
    5906, 
    4326, 
    4112, 
    6135, 
    5906, 
    4112, 
    3780, 
    3498, 
    5906, 
    6393, 
    6441, 
    6260, 
    5754, 
    4522, 
    4326, 
    5906, 
    5754, 
    4326, 
    3498, 
    3179, 
    5754, 
    6001, 
    6115, 
    5890, 
    4575, 
    4291, 
    4498, 
    5722, 
    5487, 
    5824, 
    3780, 
    4042, 
    3219, 
    6465, 
    5735, 
    5559, 
    5804, 
    6474, 
    5938, 
    4964, 
    5735, 
    6465, 
    2512, 
    2804, 
    4833, 
    3292, 
    4781, 
    2952, 
    4010, 
    4147, 
    4360, 
    3245, 
    4427, 
    2904, 
    5979, 
    6355, 
    5841, 
    4575, 
    4750, 
    6486, 
    4291, 
    4575, 
    2828, 
    4498, 
    4674, 
    4750, 
    2528, 
    2952, 
    1912, 
    5022, 
    4955, 
    2932, 
    3274, 
    5022, 
    2932, 
    4872, 
    3897, 
    5022, 
    2956, 
    4964, 
    2591, 
    2956, 
    4723, 
    4964, 
    6538, 
    5483, 
    5829, 
    5735, 
    6457, 
    5559, 
    5676, 
    5483, 
    6411, 
    5559, 
    6457, 
    6411, 
    4636, 
    4450, 
    5676, 
    4239, 
    6232, 
    5984, 
    6249, 
    5581, 
    5651, 
    5683, 
    6459, 
    5829, 
    5904, 
    5581, 
    6249, 
    5493, 
    6028, 
    6459, 
    5765, 
    5617, 
    5904, 
    5779, 
    5617, 
    5765, 
    5470, 
    5779, 
    5602, 
    5470, 
    5724, 
    5779, 
    6416, 
    6512, 
    5509, 
    6462, 
    5841, 
    5695, 
    6338, 
    5979, 
    6275, 
    6208, 
    6089, 
    5617, 
    5779, 
    6208, 
    5617, 
    5546, 
    6558, 
    6208, 
    6558, 
    6426, 
    6452, 
    6519, 
    6349, 
    5657, 
    6475, 
    6519, 
    5657, 
    6562, 
    6464, 
    6293, 
    6426, 
    6562, 
    6519, 
    6426, 
    6464, 
    6562, 
    6452, 
    6426, 
    6519, 
    6364, 
    6476, 
    6353, 
    6354, 
    6558, 
    6452, 
    5546, 
    5724, 
    6426, 
    6375, 
    6481, 
    5945, 
    6476, 
    6354, 
    6452, 
    6559, 
    6476, 
    6364, 
    6543, 
    6559, 
    6364, 
    6539, 
    6476, 
    6559, 
    6355, 
    6354, 
    6476, 
    5841, 
    6355, 
    6482, 
    6476, 
    6452, 
    6353, 
    5979, 
    6354, 
    6355, 
    5979, 
    6089, 
    6354, 
    6558, 
    6089, 
    6208, 
    6426, 
    6558, 
    5546, 
    6354, 
    6089, 
    6558, 
    5790, 
    2478, 
    5628, 
    2558, 
    5981, 
    5790, 
    2702, 
    2724, 
    3096, 
    3407, 
    4539, 
    4708, 
    3309, 
    2550, 
    2955, 
    3118, 
    3309, 
    2969, 
    3445, 
    6174, 
    4132, 
    3118, 
    3445, 
    3309, 
    3118, 
    3982, 
    3445, 
    4799, 
    4953, 
    3424, 
    2724, 
    4438, 
    3600, 
    5887, 
    2724, 
    2702, 
    3078, 
    5887, 
    2702, 
    3078, 
    4708, 
    5887, 
    3616, 
    2550, 
    3309, 
    3096, 
    3869, 
    3424, 
    3600, 
    2591, 
    4351, 
    2724, 
    3600, 
    3096, 
    6434, 
    5583, 
    2550, 
    3885, 
    6434, 
    3616, 
    6564, 
    4140, 
    5804, 
    6434, 
    6564, 
    6549, 
    3885, 
    4140, 
    6564, 
    4132, 
    3885, 
    3616, 
    3445, 
    4132, 
    3616, 
    3424, 
    3869, 
    4132, 
    5810, 
    6475, 
    5657, 
    6467, 
    6465, 
    5559, 
    5979, 
    6338, 
    6089, 
    5651, 
    5581, 
    5748, 
    6411, 
    5651, 
    5559, 
    5829, 
    5705, 
    5518, 
    6459, 
    6249, 
    5829, 
    5493, 
    6459, 
    5683, 
    5904, 
    6249, 
    6459, 
    6538, 
    6411, 
    5483, 
    5651, 
    6538, 
    5829, 
    5651, 
    6411, 
    6538, 
    5602, 
    6028, 
    3265, 
    3869, 
    4140, 
    3885, 
    3845, 
    5470, 
    3573, 
    3600, 
    4351, 
    4140, 
    4636, 
    2552, 
    3629, 
    3629, 
    4450, 
    4636, 
    2702, 
    3096, 
    4953, 
    6496, 
    965, 
    1749, 
    6496, 
    5821, 
    965, 
    3003, 
    6095, 
    2616, 
    3003, 
    3340, 
    6390, 
    6298, 
    5369, 
    684, 
    5480, 
    6298, 
    5821, 
    5480, 
    6306, 
    6298, 
    1294, 
    5964, 
    1039, 
    5335, 
    3587, 
    3281, 
    5848, 
    5588, 
    6437, 
    5579, 
    5753, 
    5238, 
    5579, 
    6326, 
    5753, 
    6368, 
    5643, 
    5678, 
    3587, 
    6368, 
    2582, 
    5848, 
    5643, 
    6368, 
    5753, 
    5848, 
    5335, 
    5753, 
    5588, 
    5848, 
    3299, 
    2757, 
    2534, 
    3281, 
    3605, 
    2940, 
    3688, 
    2702, 
    2894, 
    3605, 
    5969, 
    5774, 
    3078, 
    2702, 
    3688, 
    4047, 
    4028, 
    1933, 
    673, 
    4047, 
    1933, 
    3083, 
    2707, 
    4271, 
    5323, 
    4645, 
    4821, 
    5628, 
    5271, 
    5371, 
    5097, 
    5376, 
    5226, 
    2940, 
    3299, 
    2534, 
    5981, 
    3688, 
    5790, 
    3299, 
    5981, 
    2757, 
    3299, 
    5774, 
    5981, 
    2779, 
    4803, 
    2238, 
    2478, 
    2679, 
    5628, 
    3309, 
    3445, 
    3616, 
    2752, 
    3118, 
    2969, 
    4222, 
    2747, 
    3994, 
    3118, 
    4211, 
    3982, 
    2752, 
    2747, 
    4211, 
    1005, 
    4794, 
    2112, 
    4803, 
    4890, 
    1686, 
    4028, 
    5452, 
    2779, 
    4890, 
    880, 
    1686, 
    4957, 
    5038, 
    4803, 
    5084, 
    3994, 
    4944, 
    1912, 
    1433, 
    2418, 
    2378, 
    1912, 
    1193, 
    1433, 
    2072, 
    2418, 
    4467, 
    2574, 
    3598, 
    5036, 
    4467, 
    4259, 
    4035, 
    5172, 
    4259, 
    3114, 
    4885, 
    5036, 
    4885, 
    2752, 
    2574, 
    5036, 
    4885, 
    4467, 
    3114, 
    2747, 
    4885, 
    1272, 
    4987, 
    5374, 
    2788, 
    798, 
    1627, 
    2196, 
    4244, 
    1627, 
    777, 
    1611, 
    2788, 
    3107, 
    2739, 
    4790, 
    4534, 
    4335, 
    4339, 
    4129, 
    4534, 
    4339, 
    5930, 
    2515, 
    3990, 
    3438, 
    5930, 
    4534, 
    3438, 
    2515, 
    5930, 
    4129, 
    4339, 
    3637, 
    5619, 
    2579, 
    4252, 
    5411, 
    4315, 
    4514, 
    2494, 
    5411, 
    4514, 
    2396, 
    1468, 
    5411, 
    1468, 
    2096, 
    4315, 
    4625, 
    1750, 
    2289, 
    6127, 
    5446, 
    2494, 
    4099, 
    1383, 
    3833, 
    6500, 
    2908, 
    3250, 
    3986, 
    6127, 
    3721, 
    3986, 
    5446, 
    6127, 
    2730, 
    2347, 
    1383, 
    6319, 
    3430, 
    1482, 
    2197, 
    6319, 
    1058, 
    3721, 
    3430, 
    6319, 
    5162, 
    3721, 
    6319, 
    1149, 
    5162, 
    2197, 
    3986, 
    3721, 
    5162, 
    1886, 
    3986, 
    1149, 
    1886, 
    5446, 
    3986, 
    6500, 
    3250, 
    4704, 
    2178, 
    1115, 
    3389, 
    5088, 
    4946, 
    5092, 
    764, 
    5088, 
    4951, 
    3075, 
    4946, 
    5088, 
    1295, 
    4443, 
    1985, 
    4229, 
    3288, 
    2948, 
    764, 
    1600, 
    5088, 
    4442, 
    3288, 
    4229, 
    4951, 
    5088, 
    5092, 
    1985, 
    4951, 
    4229, 
    1985, 
    764, 
    4951, 
    5989, 
    3594, 
    3288, 
    4630, 
    5989, 
    4442, 
    4630, 
    3594, 
    5989, 
    5092, 
    4630, 
    4442, 
    2739, 
    3107, 
    6183, 
    1985, 
    4229, 
    1295, 
    2911, 
    3438, 
    5594, 
    5542, 
    5885, 
    4881, 
    6157, 
    5913, 
    5526, 
    5054, 
    6157, 
    5186, 
    5680, 
    5913, 
    6157, 
    4909, 
    5680, 
    5054, 
    2693, 
    3069, 
    5913, 
    6125, 
    3402, 
    5592, 
    5756, 
    6125, 
    5592, 
    5913, 
    3069, 
    6125, 
    5457, 
    2992, 
    5381, 
    3154, 
    3637, 
    2798, 
    4335, 
    4534, 
    5930, 
    6183, 
    3594, 
    4630, 
    6183, 
    3864, 
    3594, 
    2739, 
    6183, 
    4630, 
    4706, 
    3864, 
    6183, 
    4534, 
    4706, 
    3438, 
    4129, 
    3864, 
    4706, 
    5930, 
    3990, 
    4335, 
    3637, 
    3905, 
    4129, 
    3905, 
    3154, 
    3473, 
    4129, 
    3905, 
    3864, 
    3637, 
    3154, 
    3905, 
    2798, 
    3637, 
    3330, 
    6342, 
    3473, 
    3761, 
    3594, 
    6342, 
    4220, 
    3905, 
    3473, 
    6342, 
    5594, 
    2497, 
    2911, 
    3107, 
    5594, 
    3438, 
    3107, 
    4790, 
    5594, 
    4126, 
    2926, 
    3267, 
    4335, 
    3990, 
    4126, 
    5951, 
    4881, 
    6502, 
    4534, 
    4129, 
    4706, 
    4538, 
    4339, 
    4335, 
    6184, 
    4538, 
    4335, 
    4126, 
    6184, 
    4335, 
    4126, 
    5951, 
    6184, 
    2992, 
    3330, 
    4538, 
    3330, 
    3637, 
    4339, 
    2515, 
    2926, 
    3990, 
    4031, 
    745, 
    1972, 
    1750, 
    4031, 
    2289, 
    1750, 
    966, 
    5120, 
    4831, 
    5120, 
    966, 
    4443, 
    1972, 
    1273, 
    2289, 
    4443, 
    1295, 
    4031, 
    1972, 
    4443, 
    4443, 
    1273, 
    4515, 
    2289, 
    4031, 
    4443, 
    4823, 
    3946, 
    2021, 
    5467, 
    4976, 
    4823, 
    3510, 
    5467, 
    2845, 
    1972, 
    4976, 
    5467, 
    1972, 
    745, 
    4976, 
    5274, 
    1952, 
    3127, 
    1698, 
    898, 
    1245, 
    2259, 
    1698, 
    1245, 
    5274, 
    3832, 
    1245, 
    1952, 
    5274, 
    1245, 
    2763, 
    3832, 
    5274, 
    1708, 
    2250, 
    2259, 
    3832, 
    2241, 
    3488, 
    1245, 
    3832, 
    2259, 
    1691, 
    2241, 
    3832, 
    914, 
    1235, 
    1708, 
    1526, 
    2683, 
    665, 
    1945, 
    1235, 
    914, 
    3061, 
    3225, 
    3393, 
    2681, 
    3061, 
    2700, 
    2876, 
    872, 
    3981, 
    2038, 
    2876, 
    2681, 
    3714, 
    2972, 
    3419, 
    2876, 
    3981, 
    3225, 
    2578, 
    2972, 
    3714, 
    2235, 
    2578, 
    1681, 
    3814, 
    3093, 
    4076, 
    3814, 
    3537, 
    3419, 
    3405, 
    3690, 
    2529, 
    3393, 
    3537, 
    3690, 
    2876, 
    3225, 
    3061, 
    4076, 
    3093, 
    2718, 
    3690, 
    3814, 
    5770, 
    3690, 
    3537, 
    3814, 
    3225, 
    3537, 
    3393, 
    3419, 
    3093, 
    3814, 
    3714, 
    3419, 
    3537, 
    2972, 
    3312, 
    3419, 
    6233, 
    3308, 
    2968, 
    6097, 
    6233, 
    2968, 
    3619, 
    3312, 
    6233, 
    3419, 
    3312, 
    3093, 
    2972, 
    4898, 
    6505, 
    3537, 
    3225, 
    3714, 
    5749, 
    3076, 
    5805, 
    3405, 
    5749, 
    3690, 
    3405, 
    3076, 
    5749, 
    5805, 
    3061, 
    3393, 
    5749, 
    5805, 
    3393, 
    3076, 
    2700, 
    5805, 
    5043, 
    3884, 
    4898, 
    2235, 
    5043, 
    2578, 
    2235, 
    1213, 
    5043, 
    3312, 
    3619, 
    3093, 
    4208, 
    4292, 
    5263, 
    2139, 
    4208, 
    1547, 
    4208, 
    4404, 
    4292, 
    3619, 
    3888, 
    2718, 
    4142, 
    1945, 
    694, 
    2573, 
    4139, 
    3888, 
    4817, 
    4062, 
    2250, 
    2573, 
    4817, 
    4139, 
    2573, 
    4971, 
    4817, 
    3912, 
    4160, 
    2612, 
    5263, 
    694, 
    1547, 
    4139, 
    4142, 
    3888, 
    4139, 
    1945, 
    4142, 
    5263, 
    4142, 
    694, 
    4208, 
    5263, 
    1547, 
    5161, 
    4142, 
    5263, 
    2718, 
    5161, 
    4292, 
    3888, 
    4142, 
    5161, 
    3642, 
    4566, 
    2123, 
    4817, 
    2250, 
    1235, 
    3912, 
    4062, 
    3801, 
    3912, 
    1698, 
    4062, 
    2439, 
    665, 
    2683, 
    2123, 
    795, 
    1024, 
    1185, 
    4509, 
    4814, 
    4307, 
    4509, 
    3922, 
    16, 
    2218, 
    17, 
    4859, 
    1051, 
    1185, 
    2218, 
    4859, 
    1185, 
    1658, 
    843, 
    5157, 
    3738, 
    2816, 
    3450, 
    4380, 
    1970, 
    1268, 
    5388, 
    739, 
    1970, 
    5926, 
    5388, 
    1970, 
    4380, 
    5926, 
    1970, 
    4380, 
    1498, 
    5926, 
    699, 
    1000, 
    5388, 
    4484, 
    1489, 
    3577, 
    4050, 
    2107, 
    4484, 
    1949, 
    4050, 
    707, 
    990, 
    2107, 
    4050, 
    4697, 
    990, 
    4110, 
    6116, 
    4697, 
    4324, 
    4524, 
    2519, 
    5320, 
    32, 
    6672, 
    33, 
    2255, 
    6672, 
    31, 
    6672, 
    2255, 
    34, 
    33, 
    6672, 
    34, 
    32, 
    31, 
    6672, 
    2255, 
    35, 
    34, 
    4963, 
    1843, 
    2814, 
    358, 
    664, 
    359, 
    2058, 
    703, 
    1409, 
    2745, 
    1352, 
    908, 
    364, 
    5550, 
    908, 
    3346, 
    2122, 
    3229, 
    3229, 
    2122, 
    1525, 
    2832, 
    3182, 
    5064, 
    3539, 
    3650, 
    3346, 
    361, 
    1023, 
    362, 
    2122, 
    360, 
    1525, 
    3958, 
    664, 
    2634, 
    3920, 
    2745, 
    3650, 
    2122, 
    361, 
    360, 
    3958, 
    3229, 
    1525, 
    664, 
    3958, 
    1525, 
    3021, 
    4405, 
    3958, 
    1023, 
    361, 
    2122, 
    359, 
    1525, 
    360, 
    664, 
    1525, 
    359, 
    820, 
    1884, 
    639, 
    356, 
    820, 
    639, 
    4678, 
    355, 
    638, 
    2207, 
    4678, 
    638, 
    2207, 
    1646, 
    4678, 
    638, 
    354, 
    1164, 
    2730, 
    354, 
    353, 
    637, 
    2730, 
    353, 
    1383, 
    1164, 
    2730, 
    637, 
    2347, 
    2730, 
    871, 
    2207, 
    1164, 
    1842, 
    4931, 
    5211, 
    6241, 
    1381, 
    4299, 
    4731, 
    6241, 
    4299, 
    4841, 
    1903, 
    6241, 
    2948, 
    4625, 
    2289, 
    6342, 
    3864, 
    3905, 
    4434, 
    4220, 
    3761, 
    4252, 
    4625, 
    4026, 
    3288, 
    4220, 
    4434, 
    5457, 
    5570, 
    5709, 
    5732, 
    5556, 
    5718, 
    3473, 
    5732, 
    5718, 
    5562, 
    5738, 
    5732, 
    2798, 
    5562, 
    3154, 
    5738, 
    5556, 
    5732, 
    5709, 
    6516, 
    5562, 
    6372, 
    5883, 
    6013, 
    6420, 
    6372, 
    6371, 
    6215, 
    6420, 
    6371, 
    6516, 
    5527, 
    6420, 
    5738, 
    6516, 
    6420, 
    5738, 
    5562, 
    6516, 
    5527, 
    5883, 
    6372, 
    6518, 
    5794, 
    5420, 
    6518, 
    4026, 
    3761, 
    2579, 
    5619, 
    5420, 
    4252, 
    4026, 
    5619, 
    966, 
    4252, 
    2579, 
    966, 
    1750, 
    4252, 
    4625, 
    2948, 
    4434, 
    4026, 
    4625, 
    4434, 
    4252, 
    1750, 
    4625, 
    3288, 
    3594, 
    4220, 
    4706, 
    3107, 
    3438, 
    6342, 
    3594, 
    3864, 
    3761, 
    4220, 
    6342, 
    3761, 
    4026, 
    4434, 
    3288, 
    4442, 
    5989, 
    1295, 
    4229, 
    2948, 
    6183, 
    3107, 
    4706, 
    5877, 
    5381, 
    5284, 
    5756, 
    5877, 
    5526, 
    6431, 
    5570, 
    5457, 
    5533, 
    6431, 
    5877, 
    5533, 
    5570, 
    6431, 
    6395, 
    4196, 
    4314, 
    2798, 
    3330, 
    5457, 
    5168, 
    5580, 
    5591, 
    3820, 
    868, 
    2886, 
    4299, 
    5830, 
    3543, 
    5684, 
    868, 
    3820, 
    5830, 
    5684, 
    3820, 
    3543, 
    5830, 
    3820, 
    4299, 
    1381, 
    5830, 
    1491, 
    5591, 
    5684, 
    4678, 
    356, 
    355, 
    1680, 
    1646, 
    2207, 
    6229, 
    6013, 
    6312, 
    6395, 
    6013, 
    6229, 
    5537, 
    6126, 
    4314, 
    5537, 
    5716, 
    6550, 
    6550, 
    5716, 
    6463, 
    871, 
    4099, 
    4462, 
    4354, 
    5794, 
    6016, 
    3833, 
    3620, 
    3313, 
    4099, 
    3833, 
    3313, 
    4462, 
    4099, 
    3313, 
    1164, 
    1383, 
    4099, 
    1383, 
    4875, 
    3833, 
    3560, 
    3250, 
    3889, 
    4143, 
    3250, 
    2908, 
    6372, 
    6420, 
    5527, 
    6420, 
    5878, 
    5738, 
    6557, 
    3620, 
    6301, 
    5716, 
    6557, 
    6463, 
    3313, 
    3620, 
    6557, 
    5898, 
    5878, 
    6215, 
    4143, 
    5898, 
    3889, 
    6016, 
    5794, 
    5540, 
    4143, 
    6016, 
    5898, 
    4143, 
    4354, 
    6016, 
    5556, 
    5738, 
    5878, 
    5898, 
    6016, 
    5878, 
    5540, 
    5718, 
    5556, 
    3620, 
    3560, 
    3889, 
    3833, 
    3560, 
    3620, 
    1383, 
    2347, 
    4875, 
    5556, 
    5878, 
    6016, 
    3250, 
    4143, 
    3889, 
    2908, 
    2494, 
    4354, 
    4704, 
    4875, 
    3430, 
    5718, 
    3761, 
    3473, 
    3154, 
    5732, 
    3473, 
    5540, 
    6518, 
    5718, 
    3154, 
    5562, 
    5732, 
    5794, 
    4514, 
    5420, 
    5556, 
    6016, 
    5540, 
    4354, 
    4514, 
    5794, 
    2908, 
    4354, 
    4143, 
    5420, 
    4315, 
    2579, 
    6518, 
    5540, 
    5794, 
    4026, 
    6518, 
    5619, 
    3761, 
    5718, 
    6518, 
    4514, 
    4315, 
    5420, 
    2494, 
    4514, 
    4354, 
    2494, 
    5446, 
    5411, 
    2234, 
    820, 
    1646, 
    871, 
    1164, 
    4099, 
    1212, 
    820, 
    2234, 
    820, 
    356, 
    1646, 
    358, 
    357, 
    1884, 
    2207, 
    638, 
    1164, 
    1680, 
    2207, 
    871, 
    1646, 
    356, 
    4678, 
    1482, 
    637, 
    636, 
    6500, 
    3721, 
    6127, 
    2908, 
    6500, 
    6127, 
    4704, 
    3721, 
    6500, 
    2347, 
    637, 
    1482, 
    1058, 
    352, 
    351, 
    1058, 
    636, 
    352, 
    2197, 
    351, 
    1074, 
    5905, 
    2197, 
    1074, 
    1149, 
    3986, 
    5162, 
    1164, 
    354, 
    2730, 
    1482, 
    636, 
    1058, 
    5905, 
    1410, 
    5443, 
    5550, 
    363, 
    1023, 
    908, 
    5550, 
    2745, 
    364, 
    363, 
    5550, 
    1884, 
    820, 
    1212, 
    1928, 
    1884, 
    1212, 
    357, 
    639, 
    1884, 
    5211, 
    4931, 
    1055, 
    5430, 
    5346, 
    5211, 
    1177, 
    5430, 
    1055, 
    1177, 
    4841, 
    5430, 
    1092, 
    1842, 
    5211, 
    3346, 
    1023, 
    2122, 
    3539, 
    3346, 
    3229, 
    3958, 
    4405, 
    3229, 
    3650, 
    2745, 
    3346, 
    3394, 
    3650, 
    3539, 
    3394, 
    3063, 
    3920, 
    2745, 
    1023, 
    3346, 
    5203, 
    5075, 
    5178, 
    4765, 
    2859, 
    2233, 
    3140, 
    4765, 
    1209, 
    3140, 
    2781, 
    4765, 
    1729, 
    4941, 
    5203, 
    4941, 
    2275, 
    2887, 
    2233, 
    1679, 
    1773, 
    5990, 
    2781, 
    5453, 
    2859, 
    5990, 
    2438, 
    4765, 
    2781, 
    5990, 
    1926, 
    3140, 
    1209, 
    1926, 
    2430, 
    3892, 
    2859, 
    1679, 
    2233, 
    1209, 
    4765, 
    2233, 
    2438, 
    2470, 
    2886, 
    868, 
    992, 
    1679, 
    2943, 
    1773, 
    992, 
    5591, 
    1491, 
    5168, 
    992, 
    5591, 
    5580, 
    868, 
    5684, 
    5591, 
    2538, 
    3095, 
    2943, 
    1209, 
    2309, 
    1320, 
    2233, 
    1773, 
    2309, 
    834, 
    3063, 
    4752, 
    2948, 
    3288, 
    4434, 
    5680, 
    6157, 
    5054, 
    5709, 
    5527, 
    6516, 
    2798, 
    5709, 
    5562, 
    5570, 
    5527, 
    5709, 
    5381, 
    6431, 
    5457, 
    5533, 
    5527, 
    5570, 
    5913, 
    6125, 
    5756, 
    6395, 
    3964, 
    4196, 
    6013, 
    6395, 
    6126, 
    6229, 
    3964, 
    6395, 
    5883, 
    6312, 
    6013, 
    5592, 
    3698, 
    6229, 
    6130, 
    2992, 
    2602, 
    5885, 
    6130, 
    2602, 
    5381, 
    2992, 
    6130, 
    5526, 
    5877, 
    5284, 
    5186, 
    5526, 
    5284, 
    6229, 
    3698, 
    3964, 
    6312, 
    5592, 
    6229, 
    5533, 
    6312, 
    5883, 
    5756, 
    5592, 
    6312, 
    5877, 
    5756, 
    5533, 
    5526, 
    5913, 
    5756, 
    3402, 
    3698, 
    5592, 
    5457, 
    3330, 
    2992, 
    5420, 
    5619, 
    6518, 
    5988, 
    1381, 
    1903, 
    4909, 
    5988, 
    1903, 
    4909, 
    5860, 
    6384, 
    3233, 
    1971, 
    744, 
    3543, 
    3233, 
    4299, 
    1491, 
    5684, 
    1381, 
    3820, 
    2886, 
    2470, 
    5081, 
    2887, 
    1272, 
    3543, 
    5081, 
    3233, 
    3543, 
    2470, 
    5081, 
    6241, 
    4731, 
    4994, 
    1320, 
    2001, 
    1926, 
    2233, 
    2309, 
    1209, 
    5353, 
    4356, 
    4552, 
    2475, 
    5353, 
    4778, 
    5258, 
    4356, 
    5353, 
    4200, 
    5258, 
    2891, 
    4145, 
    4356, 
    5258, 
    5796, 
    2515, 
    2891, 
    2475, 
    5796, 
    2891, 
    2926, 
    2515, 
    5796, 
    3421, 
    3095, 
    2538, 
    3836, 
    3421, 
    3267, 
    4318, 
    3056, 
    1320, 
    3421, 
    4318, 
    3095, 
    4102, 
    3056, 
    4318, 
    3267, 
    3862, 
    4126, 
    6423, 
    4881, 
    5951, 
    2943, 
    5532, 
    2538, 
    5033, 
    4881, 
    6423, 
    992, 
    868, 
    5591, 
    5860, 
    4909, 
    5054, 
    5532, 
    5580, 
    5033, 
    6384, 
    1381, 
    5988, 
    5358, 
    1903, 
    1177, 
    5680, 
    4909, 
    5358, 
    6157, 
    5526, 
    5186, 
    2693, 
    5913, 
    5680, 
    3069, 
    3402, 
    6125, 
    5542, 
    4881, 
    5033, 
    5168, 
    5860, 
    5033, 
    5186, 
    5284, 
    5885, 
    5860, 
    5542, 
    5033, 
    1491, 
    1381, 
    6384, 
    5054, 
    5542, 
    5860, 
    4229, 
    4951, 
    4442, 
    3969, 
    2497, 
    3702, 
    4855, 
    3969, 
    3702, 
    5758, 
    3891, 
    6332, 
    2515, 
    2911, 
    2891, 
    2515, 
    3438, 
    2911, 
    4102, 
    2676, 
    3056, 
    3836, 
    4102, 
    3421, 
    3836, 
    4778, 
    4102, 
    2926, 
    3836, 
    3267, 
    2475, 
    2891, 
    5353, 
    6384, 
    5860, 
    5168, 
    1491, 
    6384, 
    5168, 
    5988, 
    4909, 
    6384, 
    6502, 
    6184, 
    5951, 
    2992, 
    6502, 
    2602, 
    4538, 
    6184, 
    6502, 
    5580, 
    2943, 
    992, 
    5033, 
    5580, 
    5168, 
    5532, 
    2943, 
    5580, 
    3075, 
    5088, 
    1600, 
    3969, 
    4200, 
    2911, 
    2458, 
    3891, 
    3623, 
    4200, 
    2891, 
    2911, 
    5758, 
    4200, 
    3969, 
    6332, 
    5258, 
    4200, 
    5758, 
    6332, 
    4200, 
    4145, 
    5258, 
    6332, 
    2458, 
    4145, 
    3891, 
    2875, 
    3224, 
    4145, 
    3095, 
    1773, 
    2943, 
    1794, 
    1025, 
    1863, 
    1579, 
    2164, 
    3390, 
    4963, 
    4395, 
    1093, 
    4116, 
    5385, 
    5461, 
    5102, 
    4395, 
    4963, 
    3057, 
    4595, 
    1794, 
    3057, 
    3390, 
    4595, 
    1980, 
    759, 
    1174, 
    2212, 
    1980, 
    1174, 
    4653, 
    2286, 
    2598, 
    2989, 
    4653, 
    2598, 
    4470, 
    5160, 
    5185, 
    2286, 
    1289, 
    1652, 
    830, 
    2441, 
    1652, 
    1744, 
    958, 
    3574, 
    958, 
    1744, 
    830, 
    2155, 
    3489, 
    4152, 
    1567, 
    2155, 
    4152, 
    4355, 
    2580, 
    4144, 
    4727, 
    4662, 
    4900, 
    5869, 
    4662, 
    4551, 
    4355, 
    6479, 
    4551, 
    3740, 
    4662, 
    5869, 
    3451, 
    4486, 
    4662, 
    4628, 
    2925, 
    2514, 
    4628, 
    4439, 
    2925, 
    2580, 
    5421, 
    4114, 
    4551, 
    4439, 
    4628, 
    5831, 
    6479, 
    4355, 
    3740, 
    3451, 
    4662, 
    4225, 
    3266, 
    4439, 
    958, 
    3314, 
    3574, 
    4144, 
    2973, 
    3890, 
    5456, 
    2795, 
    2990, 
    5640, 
    5340, 
    3773, 
    4263, 
    5640, 
    4037, 
    2514, 
    5340, 
    5640, 
    3489, 
    2795, 
    3773, 
    5340, 
    3489, 
    3773, 
    3266, 
    4152, 
    2925, 
    3266, 
    1567, 
    4152, 
    2155, 
    1078, 
    3489, 
    1432, 
    2924, 
    6383, 
    1377, 
    1031, 
    18, 
    3819, 
    1281, 
    1377, 
    3877, 
    4172, 
    940, 
    3877, 
    2734, 
    3104, 
    3025, 
    1876, 
    3300, 
    3877, 
    3104, 
    3433, 
    4172, 
    3877, 
    2639, 
    2959, 
    4172, 
    2639, 
    2080, 
    940, 
    4172, 
    940, 
    1725, 
    3877, 
    2564, 
    1139, 
    3025, 
    1444, 
    1281, 
    2080, 
    26, 
    591, 
    1281, 
    5910, 
    2374, 
    1429, 
    989, 
    5910, 
    2713, 
    4457, 
    2374, 
    5910, 
    3851, 
    4457, 
    2106, 
    1855, 
    2374, 
    4457, 
    2175, 
    3618, 
    1108, 
    4457, 
    989, 
    2106, 
    5361, 
    3189, 
    3786, 
    4788, 
    5361, 
    4420, 
    4788, 
    3505, 
    5361, 
    1108, 
    3618, 
    3627, 
    3980, 
    1693, 
    2246, 
    4788, 
    4420, 
    3980, 
    1230, 
    4788, 
    2246, 
    3505, 
    3189, 
    5361, 
    2982, 
    3320, 
    3980, 
    3627, 
    6071, 
    2589, 
    3320, 
    893, 
    1693, 
    6071, 
    6182, 
    2982, 
    2577, 
    893, 
    3320, 
    4739, 
    2307, 
    1771, 
    2070, 
    4739, 
    2713, 
    2070, 
    925, 
    4739, 
    3596, 
    2554, 
    2526, 
    2070, 
    3596, 
    925, 
    2839, 
    3189, 
    3596, 
    2374, 
    3092, 
    4619, 
    3505, 
    1940, 
    2953, 
    925, 
    3866, 
    4739, 
    6041, 
    1254, 
    4058, 
    2526, 
    2264, 
    1716, 
    3023, 
    6138, 
    2636, 
    4991, 
    3433, 
    3104, 
    6555, 
    5577, 
    5541, 
    6438, 
    6555, 
    5541, 
    6425, 
    6439, 
    6555, 
    3493, 
    5746, 
    3777, 
    3493, 
    5577, 
    5746, 
    6341, 
    5073, 
    4934, 
    6444, 
    6341, 
    5968, 
    5347, 
    6444, 
    5968, 
    5625, 
    6341, 
    6444, 
    5625, 
    5948, 
    6361, 
    5661, 
    5401, 
    5071, 
    6360, 
    5661, 
    5071, 
    6361, 
    5813, 
    6360, 
    5073, 
    6361, 
    6360, 
    6341, 
    5625, 
    6361, 
    5614, 
    5948, 
    5625, 
    6438, 
    5541, 
    6313, 
    6438, 
    6425, 
    6555, 
    6236, 
    6545, 
    6313, 
    6381, 
    6425, 
    6438, 
    5614, 
    4991, 
    6439, 
    6381, 
    5614, 
    6425, 
    6454, 
    6236, 
    5558, 
    5813, 
    6454, 
    5661, 
    5813, 
    6381, 
    6545, 
    4933, 
    4761, 
    5073, 
    5431, 
    4214, 
    5347, 
    4473, 
    3025, 
    3723, 
    4908, 
    2150, 
    3951, 
    723, 
    4635, 
    1563, 
    3951, 
    1139, 
    2190, 
    4908, 
    3951, 
    2190, 
    2150, 
    1072, 
    3951, 
    1335, 
    3455, 
    3941, 
    815, 
    2715, 
    2011, 
    3134, 
    1640, 
    4039, 
    3090, 
    3134, 
    2772, 
    815, 
    1640, 
    3134, 
    2713, 
    1771, 
    989, 
    4457, 
    5910, 
    989, 
    1429, 
    2070, 
    2713, 
    4389, 
    1317, 
    1999, 
    790, 
    4763, 
    1999, 
    3743, 
    1771, 
    2307, 
    4998, 
    3743, 
    2632, 
    4008, 
    5112, 
    5234, 
    2713, 
    4739, 
    1771, 
    3131, 
    2715, 
    3090, 
    3038, 
    2852, 
    3370, 
    3455, 
    2715, 
    3131, 
    3370, 
    3201, 
    3671, 
    1335, 
    2011, 
    3455, 
    4571, 
    5462, 
    3008, 
    5462, 
    3450, 
    2816, 
    3008, 
    5462, 
    2621, 
    3124, 
    3450, 
    5462, 
    3914, 
    4161, 
    2759, 
    5462, 
    2816, 
    2621, 
    4161, 
    4375, 
    3124, 
    3738, 
    739, 
    1574, 
    4375, 
    4567, 
    3450, 
    4567, 
    4740, 
    3738, 
    1574, 
    2161, 
    2816, 
    1692, 
    974, 
    2098, 
    4556, 
    4903, 
    892, 
    5350, 
    1759, 
    974, 
    3514, 
    1939, 
    4848, 
    2114, 
    3514, 
    1008, 
    2114, 
    688, 
    3514, 
    5326, 
    1540, 
    5415, 
    2957, 
    5326, 
    1989, 
    688, 
    1540, 
    5326, 
    3518, 
    2480, 
    5313, 
    2436, 
    3518, 
    2137, 
    3206, 
    2480, 
    3518, 
    5496, 
    3834, 
    2856, 
    4100, 
    5496, 
    3206, 
    4100, 
    3834, 
    5496, 
    4316, 
    4100, 
    2436, 
    1047, 
    4316, 
    2436, 
    1808, 
    3551, 
    4316, 
    6269, 
    2898, 
    4862, 
    4316, 
    6269, 
    4100, 
    3239, 
    2898, 
    6269, 
    2856, 
    2896, 
    3206, 
    2436, 
    4100, 
    3206, 
    1627, 
    798, 
    2856, 
    805, 
    1545, 
    693, 
    4316, 
    1047, 
    1808, 
    798, 
    2896, 
    2856, 
    2137, 
    1047, 
    2436, 
    2006, 
    2137, 
    1545, 
    1329, 
    1047, 
    2137, 
    2006, 
    1329, 
    2137, 
    2516, 
    3258, 
    1290, 
    1632, 
    3999, 
    805, 
    3268, 
    3258, 
    2516, 
    3999, 
    5700, 
    2504, 
    2754, 
    3121, 
    3447, 
    2504, 
    2916, 
    2927, 
    4087, 
    6055, 
    1981, 
    6165, 
    4087, 
    2586, 
    2979, 
    6165, 
    2586, 
    2979, 
    1001, 
    6397, 
    4302, 
    4423, 
    6055, 
    4087, 
    1981, 
    760, 
    1290, 
    5221, 
    1981, 
    2896, 
    798, 
    2004, 
    4353, 
    5085, 
    2004, 
    2480, 
    3206, 
    2896, 
    1324, 
    4353, 
    2004, 
    1545, 
    2137, 
    3518, 
    805, 
    2006, 
    1545, 
    2749, 
    3296, 
    4637, 
    5228, 
    2824, 
    3176, 
    3603, 
    5228, 
    3296, 
    5060, 
    2824, 
    5228, 
    2395, 
    4588, 
    1466, 
    2395, 
    1883, 
    4760, 
    2555, 
    4452, 
    1670, 
    4760, 
    4783, 
    2824, 
    6030, 
    860, 
    1670, 
    4452, 
    6030, 
    1670, 
    4452, 
    5932, 
    6030, 
    3939, 
    3495, 
    3176, 
    6057, 
    4414, 
    3939, 
    4414, 
    2034, 
    3939, 
    2034, 
    860, 
    3495, 
    4783, 
    2482, 
    2898, 
    4783, 
    4760, 
    2482, 
    4613, 
    4783, 
    2898, 
    4613, 
    6057, 
    4783, 
    4588, 
    2395, 
    4760, 
    2669, 
    5435, 
    1466, 
    1883, 
    2482, 
    4760, 
    1372, 
    2110, 
    2034, 
    1778, 
    1001, 
    2342, 
    2110, 
    1499, 
    2034, 
    1001, 
    2110, 
    1372, 
    5272, 
    4713, 
    2110, 
    2586, 
    5372, 
    2979, 
    4891, 
    4713, 
    5272, 
    1109, 
    4891, 
    5372, 
    1109, 
    1856, 
    4891, 
    3779, 
    860, 
    2034, 
    1499, 
    3779, 
    2034, 
    1499, 
    2416, 
    3779, 
    4713, 
    1499, 
    2110, 
    1001, 
    5272, 
    2110, 
    5504, 
    1856, 
    3659, 
    5504, 
    4891, 
    1856, 
    3357, 
    5504, 
    3659, 
    3357, 
    4713, 
    5504, 
    2586, 
    1596, 
    2176, 
    4891, 
    5272, 
    5372, 
    1778, 
    6397, 
    1001, 
    4423, 
    2315, 
    1329, 
    6165, 
    4302, 
    4087, 
    1778, 
    2315, 
    4302, 
    6397, 
    1778, 
    4302, 
    6165, 
    6397, 
    4302, 
    6165, 
    2979, 
    6397, 
    3470, 
    1950, 
    1243, 
    1109, 
    5139, 
    1856, 
    708, 
    1950, 
    3470, 
    3700, 
    3968, 
    3183, 
    1513, 
    3700, 
    3183, 
    2675, 
    5436, 
    3700, 
    1641, 
    2204, 
    762, 
    2830, 
    4691, 
    5436, 
    2756, 
    4878, 
    2737, 
    3589, 
    2073, 
    1434, 
    2596, 
    931, 
    2073, 
    3589, 
    2596, 
    2073, 
    1869, 
    1128, 
    2596, 
    6268, 
    2312, 
    1324, 
    2386, 
    4373, 
    1869, 
    1774, 
    2312, 
    3911, 
    2510, 
    2004, 
    798, 
    2184, 
    2510, 
    1611, 
    2184, 
    3563, 
    2510, 
    2795, 
    3489, 
    1078, 
    2987, 
    1880, 
    2888, 
    2471, 
    2987, 
    2888, 
    2945, 
    2393, 
    2987, 
    3890, 
    3314, 
    3621, 
    2393, 
    1880, 
    2987, 
    4749, 
    1719, 
    931, 
    2596, 
    4749, 
    931, 
    1128, 
    2184, 
    4749, 
    4662, 
    4727, 
    4551, 
    1963, 
    4225, 
    4900, 
    4628, 
    2514, 
    4114, 
    4807, 
    2267, 
    1719, 
    4749, 
    4807, 
    1719, 
    2184, 
    1611, 
    4807, 
    1611, 
    1260, 
    2267, 
    3563, 
    2004, 
    2510, 
    777, 
    1260, 
    1611, 
    1151, 
    346, 
    345, 
    633, 
    3576, 
    3850, 
    1410, 
    346, 
    1151, 
    5385, 
    4116, 
    1437, 
    1025, 
    5385, 
    933, 
    5461, 
    2814, 
    6175, 
    5102, 
    5461, 
    5385, 
    5102, 
    4963, 
    5461, 
    4595, 
    5102, 
    1025, 
    4963, 
    2814, 
    5461, 
    1410, 
    2814, 
    2364, 
    5102, 
    5385, 
    1025, 
    6175, 
    4116, 
    5461, 
    3576, 
    1437, 
    4116, 
    5411, 
    1468, 
    4315, 
    5446, 
    2396, 
    5411, 
    2908, 
    6127, 
    2494, 
    1886, 
    2396, 
    5446, 
    2396, 
    4652, 
    2966, 
    5443, 
    2364, 
    4652, 
    2966, 
    1468, 
    2396, 
    6604, 
    343, 
    342, 
    3850, 
    6604, 
    633, 
    3850, 
    343, 
    6604, 
    4116, 
    3850, 
    3576, 
    1151, 
    343, 
    3850, 
    6205, 
    3679, 
    2966, 
    1117, 
    1263, 
    1794, 
    2197, 
    1058, 
    351, 
    5974, 
    1886, 
    1149, 
    5974, 
    4652, 
    1886, 
    5443, 
    5974, 
    1149, 
    5443, 
    4652, 
    5974, 
    6087, 
    1843, 
    6205, 
    2364, 
    6087, 
    4652, 
    2364, 
    1843, 
    6087, 
    1151, 
    6175, 
    1410, 
    4652, 
    2396, 
    1886, 
    6087, 
    2966, 
    4652, 
    6205, 
    1093, 
    3679, 
    6087, 
    6205, 
    2966, 
    1843, 
    1093, 
    6205, 
    4831, 
    966, 
    2096, 
    2164, 
    4831, 
    3679, 
    2164, 
    1579, 
    4831, 
    4395, 
    4595, 
    3390, 
    5120, 
    4031, 
    1750, 
    1579, 
    5120, 
    4831, 
    1579, 
    745, 
    5120, 
    2096, 
    966, 
    2579, 
    3679, 
    2096, 
    1468, 
    2966, 
    3679, 
    1468, 
    1093, 
    2164, 
    3679, 
    1295, 
    2948, 
    2289, 
    2347, 
    1482, 
    3430, 
    6319, 
    1482, 
    1058, 
    2197, 
    5162, 
    6319, 
    4875, 
    3560, 
    3833, 
    3430, 
    4875, 
    2347, 
    4704, 
    3560, 
    4875, 
    3721, 
    4704, 
    3430, 
    3250, 
    3560, 
    4704, 
    4315, 
    2096, 
    2579, 
    2243, 
    338, 
    337, 
    2243, 
    1227, 
    338, 
    4233, 
    4007, 
    336, 
    4233, 
    2765, 
    4007, 
    335, 
    4233, 
    336, 
    335, 
    334, 
    4233, 
    5654, 
    5957, 
    6291, 
    2213, 
    3453, 
    2765, 
    5978, 
    835, 
    993, 
    1492, 
    5635, 
    4822, 
    1492, 
    835, 
    5635, 
    4633, 
    1863, 
    933, 
    4633, 
    4810, 
    5477, 
    5978, 
    5635, 
    835, 
    2760, 
    5978, 
    3125, 
    4822, 
    5635, 
    5978, 
    6214, 
    341, 
    340, 
    339, 
    6214, 
    340, 
    3168, 
    3487, 
    6214, 
    6214, 
    1437, 
    341, 
    6450, 
    5672, 
    5477, 
    6084, 
    6450, 
    5654, 
    6084, 
    5116, 
    6450, 
    4633, 
    933, 
    3487, 
    3168, 
    4810, 
    3487, 
    2543, 
    1863, 
    4633, 
    4395, 
    5102, 
    4595, 
    3487, 
    933, 
    1437, 
    6214, 
    3487, 
    1437, 
    6389, 
    5654, 
    4007, 
    3453, 
    6389, 
    2765, 
    6084, 
    5654, 
    6389, 
    4822, 
    6084, 
    6389, 
    4975, 
    5116, 
    6084, 
    3487, 
    4810, 
    4633, 
    3168, 
    1227, 
    4961, 
    6291, 
    2243, 
    4007, 
    5654, 
    6291, 
    4007, 
    4961, 
    2243, 
    6291, 
    3168, 
    4961, 
    4810, 
    1227, 
    2243, 
    4961, 
    1117, 
    1794, 
    1863, 
    3946, 
    1355, 
    2021, 
    1263, 
    2332, 
    1794, 
    1263, 
    1355, 
    2332, 
    3679, 
    4831, 
    2096, 
    3057, 
    2332, 
    1355, 
    4182, 
    6083, 
    3946, 
    1093, 
    4395, 
    2164, 
    4595, 
    1025, 
    1794, 
    2164, 
    4395, 
    3390, 
    1093, 
    1843, 
    4963, 
    1794, 
    2332, 
    3057, 
    745, 
    4031, 
    5120, 
    3168, 
    6214, 
    339, 
    4353, 
    2312, 
    3837, 
    2788, 
    1611, 
    2510, 
    4103, 
    1234, 
    1944, 
    4490, 
    3837, 
    4282, 
    693, 
    4726, 
    1944, 
    4726, 
    5313, 
    5045, 
    4103, 
    4726, 
    4516, 
    693, 
    1545, 
    5313, 
    2312, 
    1774, 
    4282, 
    4282, 
    1774, 
    3301, 
    4490, 
    4282, 
    3607, 
    2248, 
    4490, 
    3607, 
    4103, 
    3837, 
    4490, 
    3837, 
    2312, 
    4282, 
    3563, 
    6268, 
    1324, 
    1128, 
    1869, 
    3911, 
    3607, 
    3301, 
    2562, 
    1234, 
    4490, 
    2248, 
    1234, 
    4103, 
    4490, 
    6213, 
    969, 
    3921, 
    4024, 
    5041, 
    2412, 
    896, 
    2807, 
    2053, 
    2562, 
    3301, 
    5288, 
    5041, 
    5288, 
    1494, 
    1697, 
    2562, 
    896, 
    1697, 
    2248, 
    3607, 
    996, 
    4373, 
    5330, 
    6225, 
    3204, 
    2854, 
    2053, 
    4719, 
    1403, 
    2412, 
    1904, 
    4024, 
    5040, 
    1298, 
    1082, 
    837, 
    5040, 
    1654, 
    1570, 
    1298, 
    5040, 
    2021, 
    5407, 
    837, 
    5574, 
    3302, 
    2563, 
    732, 
    6323, 
    1570, 
    6154, 
    4546, 
    4715, 
    5574, 
    6323, 
    6034, 
    6323, 
    1603, 
    6154, 
    5601, 
    1753, 
    1082, 
    2680, 
    5012, 
    5590, 
    3776, 
    3921, 
    4858, 
    4654, 
    5040, 
    1082, 
    6324, 
    1603, 
    1263, 
    5273, 
    6324, 
    1263, 
    2543, 
    5273, 
    1117, 
    5239, 
    6161, 
    5273, 
    6324, 
    6161, 
    4715, 
    1603, 
    6324, 
    4546, 
    5273, 
    6161, 
    6324, 
    4633, 
    5477, 
    6530, 
    6161, 
    4893, 
    4715, 
    5116, 
    5448, 
    5239, 
    5116, 
    2760, 
    5448, 
    5476, 
    4893, 
    2760, 
    2761, 
    5449, 
    4893, 
    5745, 
    3608, 
    3302, 
    4893, 
    5449, 
    4715, 
    2761, 
    3876, 
    5745, 
    5745, 
    5449, 
    2761, 
    5574, 
    6034, 
    3302, 
    5449, 
    6154, 
    4715, 
    3302, 
    6034, 
    5745, 
    6323, 
    732, 
    1603, 
    6034, 
    6323, 
    6154, 
    5574, 
    1570, 
    6323, 
    3615, 
    3884, 
    2439, 
    1463, 
    2235, 
    1681, 
    1463, 
    2394, 
    2235, 
    2094, 
    1463, 
    1681, 
    4624, 
    2198, 
    1152, 
    5370, 
    5319, 
    2754, 
    1632, 
    5370, 
    3999, 
    2198, 
    4624, 
    5370, 
    3793, 
    4433, 
    3167, 
    5319, 
    3121, 
    2754, 
    3793, 
    4798, 
    4433, 
    3793, 
    1463, 
    4798, 
    1745, 
    3121, 
    959, 
    1745, 
    3258, 
    3447, 
    5370, 
    1632, 
    2198, 
    5700, 
    3999, 
    2754, 
    2504, 
    805, 
    3999, 
    5370, 
    2754, 
    3999, 
    4798, 
    5319, 
    4433, 
    4798, 
    3121, 
    5319, 
    2398, 
    1697, 
    896, 
    2669, 
    2095, 
    4243, 
    5435, 
    2669, 
    979, 
    1466, 
    2095, 
    2669, 
    5435, 
    2395, 
    1466, 
    1763, 
    5435, 
    979, 
    1763, 
    5287, 
    5435, 
    2824, 
    4588, 
    4760, 
    1641, 
    762, 
    1598, 
    2405, 
    1747, 
    2288, 
    893, 
    2405, 
    1894, 
    2051, 
    1478, 
    2405, 
    1292, 
    1983, 
    1159, 
    1693, 
    1894, 
    1159, 
    4342, 
    2749, 
    2555, 
    1919, 
    4668, 
    1202, 
    4668, 
    2740, 
    4489, 
    4383, 
    844, 
    2025, 
    2877, 
    4383, 
    2025, 
    1513, 
    2425, 
    5697, 
    4668, 
    4489, 
    5867, 
    3108, 
    4668, 
    1919, 
    3108, 
    2740, 
    4668, 
    4342, 
    2228, 
    1202, 
    5060, 
    1466, 
    4588, 
    1670, 
    2228, 
    2555, 
    1670, 
    4085, 
    2228, 
    3603, 
    3293, 
    962, 
    2095, 
    3603, 
    962, 
    3296, 
    3597, 
    3603, 
    3176, 
    4637, 
    5228, 
    4217, 
    6259, 
    3991, 
    3296, 
    3867, 
    3597, 
    3867, 
    2749, 
    5867, 
    1478, 
    2101, 
    4243, 
    4637, 
    3296, 
    5228, 
    5932, 
    4637, 
    3176, 
    4452, 
    2555, 
    4637, 
    5768, 
    3779, 
    2416, 
    4085, 
    5768, 
    2416, 
    4085, 
    1670, 
    5768, 
    5697, 
    2647, 
    844, 
    1513, 
    5697, 
    4383, 
    2425, 
    2647, 
    5697, 
    5143, 
    2219, 
    3034, 
    2548, 
    4999, 
    926, 
    2647, 
    3034, 
    1659, 
    6036, 
    4677, 
    4999, 
    2219, 
    6036, 
    4999, 
    1186, 
    5158, 
    6036, 
    6000, 
    1186, 
    5143, 
    2228, 
    6000, 
    5143, 
    4085, 
    1908, 
    6000, 
    860, 
    3779, 
    5768, 
    3659, 
    1856, 
    2375, 
    1430, 
    3659, 
    2375, 
    5504, 
    4713, 
    4891, 
    5158, 
    1186, 
    1908, 
    1430, 
    4677, 
    3659, 
    1430, 
    2071, 
    4677, 
    2416, 
    1499, 
    4713, 
    4085, 
    2416, 
    1908, 
    1186, 
    6000, 
    1908, 
    1670, 
    860, 
    5768, 
    2416, 
    4713, 
    3357, 
    4325, 
    1717, 
    2265, 
    1659, 
    4325, 
    844, 
    2548, 
    1717, 
    4325, 
    2548, 
    926, 
    1717, 
    2219, 
    2548, 
    1659, 
    2219, 
    1186, 
    6036, 
    4999, 
    2071, 
    926, 
    2219, 
    4999, 
    2548, 
    4677, 
    2071, 
    4999, 
    1430, 
    3827, 
    5589, 
    1908, 
    2416, 
    3357, 
    4602, 
    6132, 
    912, 
    1430, 
    5589, 
    2071, 
    2257, 
    1706, 
    2741, 
    5589, 
    2257, 
    2741, 
    2071, 
    5589, 
    2741, 
    3827, 
    2257, 
    5589, 
    4614, 
    4415, 
    1950, 
    3508, 
    4784, 
    3789, 
    4204, 
    4415, 
    4614, 
    6277, 
    4128, 
    2061, 
    2367, 
    6277, 
    1413, 
    4014, 
    5791, 
    6277, 
    4638, 
    4968, 
    1255, 
    6277, 
    2061, 
    1413, 
    1717, 
    4128, 
    2265, 
    1717, 
    4602, 
    4128, 
    5236, 
    4950, 
    2206, 
    4456, 
    6219, 
    4640, 
    4897, 
    4950, 
    5236, 
    4559, 
    5545, 
    4736, 
    2790, 
    4559, 
    4149, 
    5545, 
    3846, 
    4736, 
    2575, 
    5545, 
    4559, 
    4113, 
    3846, 
    5545, 
    3323, 
    3632, 
    4907, 
    2559, 
    3873, 
    3900, 
    4523, 
    819, 
    1645, 
    2790, 
    3148, 
    2575, 
    2014, 
    819, 
    2970, 
    3148, 
    4558, 
    1340, 
    4736, 
    3632, 
    3900, 
    4559, 
    4736, 
    3900, 
    5863, 
    2513, 
    6287, 
    3180, 
    2675, 
    1013, 
    2324, 
    4170, 
    1787, 
    2830, 
    2675, 
    3180, 
    4345, 
    2830, 
    4170, 
    6147, 
    4134, 
    4345, 
    2575, 
    4559, 
    2790, 
    3900, 
    3873, 
    4149, 
    6168, 
    4925, 
    4511, 
    4149, 
    3873, 
    4134, 
    2575, 
    4327, 
    5545, 
    3632, 
    2559, 
    3900, 
    4310, 
    4925, 
    5062, 
    6532, 
    4431, 
    4217, 
    4609, 
    5195, 
    6532, 
    4609, 
    1983, 
    5195, 
    2985, 
    1032, 
    2128, 
    1534, 
    3757, 
    2128, 
    1340, 
    2324, 
    3322, 
    2970, 
    2575, 
    3148, 
    2958, 
    2559, 
    3632, 
    2177, 
    5062, 
    1112, 
    5062, 
    4093, 
    4310, 
    2958, 
    5062, 
    4925, 
    2177, 
    4093, 
    5062, 
    3148, 
    1340, 
    2014, 
    2970, 
    3148, 
    2014, 
    2790, 
    6147, 
    4558, 
    3352, 
    3322, 
    2324, 
    3322, 
    1032, 
    2985, 
    1787, 
    3352, 
    2324, 
    1797, 
    1032, 
    3322, 
    2985, 
    2128, 
    3757, 
    1340, 
    2985, 
    2014, 
    3899, 
    1564, 
    2151, 
    2128, 
    3899, 
    2151, 
    1032, 
    3631, 
    3899, 
    1340, 
    3322, 
    2985, 
    3352, 
    1797, 
    3322, 
    1013, 
    5009, 
    1787, 
    2336, 
    1797, 
    3352, 
    1787, 
    5009, 
    3352, 
    3226, 
    1960, 
    724, 
    1362, 
    3226, 
    2336, 
    1362, 
    4638, 
    3226, 
    1797, 
    3226, 
    724, 
    2151, 
    1073, 
    2128, 
    1032, 
    3899, 
    2128, 
    3399, 
    2714, 
    1846, 
    2167, 
    3399, 
    1096, 
    3067, 
    2714, 
    3399, 
    2151, 
    3067, 
    2688, 
    1564, 
    724, 
    3067, 
    1797, 
    3631, 
    1032, 
    724, 
    2714, 
    3067, 
    3786, 
    2839, 
    2070, 
    4619, 
    5361, 
    3786, 
    2982, 
    4420, 
    2589, 
    3980, 
    2246, 
    4788, 
    1230, 
    3505, 
    4788, 
    1230, 
    1940, 
    3505, 
    3505, 
    2953, 
    3189, 
    4009, 
    5237, 
    2770, 
    6390, 
    5321, 
    5480, 
    5821, 
    6390, 
    5480, 
    6095, 
    3003, 
    6390, 
    6298, 
    2753, 
    5369, 
    684, 
    5821, 
    6298, 
    6306, 
    5156, 
    5907, 
    3645, 
    5321, 
    3340, 
    5321, 
    5156, 
    6306, 
    2937, 
    5615, 
    2530, 
    6113, 
    5454, 
    5638, 
    5037, 
    6113, 
    3120, 
    5037, 
    2789, 
    6113, 
    6171, 
    1467, 
    684, 
    5638, 
    6171, 
    5369, 
    1226, 
    1467, 
    6171, 
    4377, 
    5425, 
    2909, 
    5425, 
    2620, 
    2495, 
    5344, 
    5425, 
    4377, 
    5344, 
    1226, 
    6171, 
    5037, 
    4886, 
    3147, 
    5454, 
    6113, 
    2789, 
    3446, 
    4886, 
    5037, 
    5907, 
    3446, 
    3120, 
    2937, 
    3278, 
    3734, 
    3343, 
    6242, 
    6402, 
    3120, 
    3446, 
    5037, 
    6286, 
    3756, 
    1029, 
    6402, 
    6286, 
    1018, 
    6402, 
    3469, 
    6286, 
    3446, 
    3734, 
    4886, 
    6286, 
    1791, 
    1018, 
    5576, 
    3998, 
    6011, 
    4886, 
    5576, 
    3469, 
    4886, 
    3734, 
    5576, 
    1029, 
    1791, 
    6286, 
    3007, 
    2495, 
    2620, 
    2789, 
    5960, 
    2620, 
    4786, 
    6139, 
    841, 
    5960, 
    3343, 
    3007, 
    2620, 
    5960, 
    3007, 
    3147, 
    3469, 
    6242, 
    1359, 
    1519, 
    6139, 
    2722, 
    2339, 
    4413, 
    3422, 
    2722, 
    1018, 
    1365, 
    2339, 
    2722, 
    4377, 
    2909, 
    1148, 
    1226, 
    5344, 
    1885, 
    5425, 
    2495, 
    2909, 
    5822, 
    6139, 
    4786, 
    5155, 
    1656, 
    1205, 
    2495, 
    4616, 
    4416, 
    6093, 
    1656, 
    5155, 
    5378, 
    6093, 
    5155, 
    4786, 
    1656, 
    6093, 
    5346, 
    1092, 
    5211, 
    6283, 
    2585, 
    5568, 
    744, 
    2978, 
    3531, 
    744, 
    1971, 
    2978, 
    3531, 
    2978, 
    2585, 
    6283, 
    3531, 
    2585, 
    3669, 
    6283, 
    3368, 
    3669, 
    3531, 
    6283, 
    1578, 
    744, 
    3531, 
    5454, 
    2789, 
    2620, 
    5344, 
    5454, 
    5425, 
    5638, 
    2753, 
    6113, 
    1148, 
    4209, 
    1885, 
    5939, 
    3396, 
    3691, 
    4789, 
    5494, 
    2685, 
    5426, 
    800, 
    2005, 
    5426, 
    3691, 
    800, 
    3396, 
    1629, 
    3691, 
    5374, 
    2978, 
    1971, 
    1272, 
    5374, 
    1971, 
    4987, 
    2776, 
    5374, 
    4290, 
    5953, 
    6521, 
    4497, 
    5646, 
    5953, 
    5524, 
    2685, 
    3065, 
    4407, 
    6309, 
    4191, 
    5876, 
    2462, 
    3227, 
    6487, 
    5876, 
    5600, 
    6010, 
    6487, 
    5600, 
    6010, 
    6309, 
    6487, 
    4407, 
    1241, 
    5876, 
    3094, 
    5923, 
    2785, 
    5923, 
    3211, 
    2861, 
    2785, 
    5923, 
    3144, 
    3094, 
    3211, 
    5923, 
    5923, 
    2861, 
    4789, 
    3524, 
    3368, 
    3211, 
    2719, 
    3803, 
    3094, 
    3803, 
    1092, 
    2163, 
    3094, 
    3803, 
    3524, 
    2719, 
    1092, 
    3803, 
    3036, 
    2861, 
    3211, 
    5568, 
    3036, 
    3368, 
    3893, 
    6026, 
    2585, 
    3893, 
    3460, 
    5481, 
    2650, 
    2861, 
    3036, 
    4767, 
    1885, 
    4209, 
    2442, 
    4767, 
    4209, 
    5646, 
    4497, 
    1467, 
    2650, 
    5646, 
    4767, 
    2650, 
    5953, 
    5646, 
    4841, 
    5346, 
    5430, 
    1680, 
    2234, 
    1646, 
    2910, 
    2846, 
    2496, 
    4258, 
    2910, 
    4034, 
    2618, 
    4258, 
    4034, 
    3005, 
    3341, 
    4466, 
    4525, 
    6533, 
    3494, 
    6531, 
    5675, 
    4137, 
    3341, 
    6531, 
    5747, 
    3341, 
    5675, 
    6531, 
    5719, 
    2823, 
    3175, 
    4137, 
    5719, 
    4349, 
    4137, 
    5020, 
    5719, 
    4648, 
    3646, 
    4272, 
    4466, 
    4648, 
    3561, 
    4466, 
    3341, 
    4648, 
    5199, 
    5131, 
    3835, 
    5395, 
    3561, 
    5131, 
    3526, 
    5395, 
    5131, 
    3214, 
    5468, 
    5395, 
    3252, 
    4466, 
    3561, 
    3511, 
    2496, 
    2445, 
    4063, 
    4283, 
    2445, 
    4051, 
    2212, 
    3162, 
    2808, 
    4051, 
    3162, 
    3791, 
    1652, 
    4051, 
    4283, 
    4491, 
    3511, 
    1652, 
    2212, 
    4051, 
    5194, 
    1488, 
    2106, 
    3609, 
    3128, 
    3452, 
    4724, 
    4617, 
    4965, 
    5106, 
    4724, 
    4965, 
    2962, 
    5106, 
    3303, 
    5194, 
    2106, 
    4548, 
    2962, 
    5194, 
    5106, 
    2962, 
    1488, 
    5194, 
    5112, 
    4008, 
    2570, 
    4548, 
    5112, 
    4724, 
    5234, 
    1771, 
    3743, 
    4548, 
    5234, 
    5112, 
    4548, 
    989, 
    5234, 
    5020, 
    4137, 
    2764, 
    5650, 
    5020, 
    3609, 
    4812, 
    2823, 
    5020, 
    5127, 
    2618, 
    4034, 
    3162, 
    5127, 
    2808, 
    3452, 
    3128, 
    5127, 
    5127, 
    3128, 
    2618, 
    5242, 
    3741, 
    3452, 
    3303, 
    3609, 
    3452, 
    5194, 
    4724, 
    5106, 
    4418, 
    2965, 
    4206, 
    2764, 
    2618, 
    3128, 
    2018, 
    958, 
    830, 
    4159, 
    1990, 
    3519, 
    1348, 
    2093, 
    2018, 
    5463, 
    2825, 
    2503, 
    3257, 
    5463, 
    2915, 
    2930, 
    2825, 
    5463, 
    1792, 
    4667, 
    3112, 
    4221, 
    4435, 
    4474, 
    2557, 
    3448, 
    3736, 
    2888, 
    1880, 
    1143, 
    2193, 
    3736, 
    1143, 
    2987, 
    3324, 
    2945, 
    2762, 
    1719, 
    2267, 
    6247, 
    3901, 
    3633, 
    5208, 
    6247, 
    4878, 
    5208, 
    4150, 
    6247, 
    5082, 
    4362, 
    5208, 
    3451, 
    4362, 
    2791, 
    3740, 
    4150, 
    4362, 
    3740, 
    4005, 
    4150, 
    3324, 
    3633, 
    2540, 
    3324, 
    2471, 
    5408, 
    5109, 
    3436, 
    2756, 
    4545, 
    4969, 
    2458, 
    3725, 
    3436, 
    4969, 
    4124, 
    3149, 
    2791, 
    4216, 
    4124, 
    3989, 
    2073, 
    931, 
    4124, 
    4333, 
    2791, 
    5082, 
    3451, 
    2791, 
    2762, 
    2267, 
    4486, 
    2762, 
    3901, 
    4005, 
    4230, 
    4545, 
    2458, 
    3623, 
    6063, 
    4712, 
    4545, 
    3317, 
    6063, 
    3623, 
    3317, 
    4712, 
    6063, 
    5270, 
    3725, 
    4969, 
    4639, 
    5270, 
    4545, 
    4639, 
    3989, 
    5270, 
    3451, 
    3740, 
    4362, 
    5109, 
    2875, 
    4969, 
    3436, 
    5109, 
    4969, 
    5845, 
    3224, 
    2875, 
    2756, 
    5845, 
    5109, 
    2756, 
    5327, 
    5845, 
    3324, 
    2540, 
    2945, 
    2471, 
    3324, 
    2987, 
    5408, 
    2737, 
    4878, 
    3324, 
    5408, 
    3633, 
    2471, 
    2737, 
    5408, 
    4551, 
    4628, 
    5421, 
    1462, 
    2330, 
    2393, 
    2393, 
    2330, 
    1792, 
    2121, 
    1143, 
    1022, 
    3728, 
    3441, 
    2963, 
    3304, 
    3728, 
    2963, 
    2930, 
    3272, 
    3728, 
    1792, 
    3112, 
    1022, 
    1792, 
    2330, 
    4667, 
    1523, 
    1623, 
    2121, 
    3947, 
    1115, 
    2178, 
    2084, 
    2583, 
    944, 
    2084, 
    1449, 
    5117, 
    4545, 
    5270, 
    4969, 
    5270, 
    3989, 
    3725, 
    3623, 
    6063, 
    4545, 
    4453, 
    4216, 
    4639, 
    1434, 
    4216, 
    4453, 
    1434, 
    2073, 
    4216, 
    4216, 
    2073, 
    4124, 
    4902, 
    2676, 
    4729, 
    3813, 
    3298, 
    2557, 
    4729, 
    3813, 
    4075, 
    4778, 
    4729, 
    2676, 
    4552, 
    3813, 
    4729, 
    3536, 
    3298, 
    3813, 
    4778, 
    5353, 
    4552, 
    3536, 
    5845, 
    5327, 
    4552, 
    4356, 
    3536, 
    3813, 
    4552, 
    3536, 
    4778, 
    3836, 
    2475, 
    4729, 
    4778, 
    4552, 
    2676, 
    4102, 
    4778, 
    2875, 
    5109, 
    5845, 
    3448, 
    2737, 
    2471, 
    4075, 
    3813, 
    2557, 
    1623, 
    4075, 
    2557, 
    794, 
    2001, 
    4902, 
    5327, 
    2737, 
    3448, 
    3536, 
    5327, 
    3298, 
    3536, 
    3224, 
    5845, 
    3149, 
    931, 
    1719, 
    4333, 
    3989, 
    4124, 
    4362, 
    5082, 
    2791, 
    3725, 
    3989, 
    4333, 
    4124, 
    931, 
    3149, 
    3149, 
    1719, 
    2762, 
    3736, 
    2888, 
    1143, 
    2557, 
    3736, 
    2193, 
    3448, 
    2888, 
    3736, 
    5327, 
    3448, 
    3298, 
    2471, 
    2888, 
    3448, 
    3298, 
    3448, 
    2557, 
    2945, 
    1462, 
    2393, 
    4878, 
    2756, 
    3436, 
    5208, 
    4878, 
    3436, 
    5082, 
    5208, 
    3436, 
    4150, 
    3901, 
    6247, 
    6247, 
    3633, 
    5408, 
    3314, 
    958, 
    2093, 
    3574, 
    2973, 
    3847, 
    1744, 
    3574, 
    2598, 
    3314, 
    2973, 
    3574, 
    1462, 
    3621, 
    2093, 
    3621, 
    2945, 
    2540, 
    2093, 
    3621, 
    3314, 
    1462, 
    2945, 
    3621, 
    3847, 
    2989, 
    2598, 
    2580, 
    3847, 
    2973, 
    2580, 
    4114, 
    3847, 
    4727, 
    4439, 
    4551, 
    4486, 
    4900, 
    4662, 
    4225, 
    4439, 
    4727, 
    5869, 
    6479, 
    3740, 
    2973, 
    4144, 
    2580, 
    3890, 
    2540, 
    4144, 
    5082, 
    3436, 
    3725, 
    4333, 
    5082, 
    3725, 
    4362, 
    4150, 
    5208, 
    4005, 
    3901, 
    4150, 
    4355, 
    4144, 
    5831, 
    4144, 
    2540, 
    4230, 
    6247, 
    5408, 
    4878, 
    2598, 
    2286, 
    1744, 
    4114, 
    3326, 
    2989, 
    5421, 
    4628, 
    4114, 
    4355, 
    5421, 
    2580, 
    4355, 
    4551, 
    5421, 
    2514, 
    3326, 
    4114, 
    4470, 
    3326, 
    4263, 
    3574, 
    3847, 
    2598, 
    3634, 
    5379, 
    5456, 
    3847, 
    4114, 
    2989, 
    2514, 
    2925, 
    5340, 
    1963, 
    728, 
    4225, 
    958, 
    2018, 
    2093, 
    1880, 
    1792, 
    1022, 
    4667, 
    2568, 
    3112, 
    4658, 
    4667, 
    2330, 
    4658, 
    4834, 
    4667, 
    4372, 
    4658, 
    1348, 
    2610, 
    4834, 
    4658, 
    4491, 
    4283, 
    4372, 
    2018, 
    4491, 
    4372, 
    830, 
    3791, 
    4491, 
    3252, 
    5468, 
    2910, 
    5286, 
    4159, 
    5189, 
    2298, 
    5286, 
    2860, 
    2298, 
    1307, 
    5286, 
    5832, 
    3802, 
    2445, 
    5468, 
    5832, 
    2846, 
    5468, 
    3214, 
    5832, 
    3992, 
    3304, 
    4221, 
    4486, 
    2267, 
    1260, 
    4900, 
    4486, 
    1260, 
    1963, 
    4900, 
    1260, 
    4225, 
    4727, 
    4900, 
    3451, 
    2762, 
    4486, 
    1348, 
    1462, 
    2093, 
    1880, 
    1022, 
    1143, 
    1348, 
    2330, 
    1462, 
    3519, 
    1990, 
    776, 
    3304, 
    5250, 
    5348, 
    5189, 
    3523, 
    3210, 
    5348, 
    5250, 
    3640, 
    3519, 
    5348, 
    3910, 
    3610, 
    3304, 
    5348, 
    3334, 
    6044, 
    5514, 
    3728, 
    3272, 
    3441, 
    2825, 
    2930, 
    2521, 
    3441, 
    3112, 
    2568, 
    2963, 
    3441, 
    2568, 
    3272, 
    3578, 
    3441, 
    5389, 
    3272, 
    2930, 
    5463, 
    5389, 
    2930, 
    3257, 
    3566, 
    5389, 
    3578, 
    1022, 
    3112, 
    2330, 
    1348, 
    4658, 
    1880, 
    2393, 
    1792, 
    1348, 
    2018, 
    4372, 
    4561, 
    1477, 
    2404, 
    4286, 
    3051, 
    3383, 
    4869, 
    5019, 
    4067, 
    1962, 
    3051, 
    4286, 
    3805, 
    1762, 
    2860, 
    3743, 
    4008, 
    5234, 
    4634, 
    3306, 
    4447, 
    5827, 
    5071, 
    5132, 
    2653, 
    3612, 
    4634, 
    6185, 
    2768, 
    3882, 
    2852, 
    3038, 
    2653, 
    2852, 
    3201, 
    3370, 
    5740, 
    2852, 
    2432, 
    4178, 
    3940, 
    2851, 
    1008, 
    4178, 
    3200, 
    3795, 
    3940, 
    4178, 
    3795, 
    3515, 
    3940, 
    2321, 
    3795, 
    1784, 
    2321, 
    3941, 
    3795, 
    3201, 
    3670, 
    3515, 
    4137, 
    5675, 
    2764, 
    4525, 
    4328, 
    4718, 
    6533, 
    4525, 
    5275, 
    5719, 
    6533, 
    4349, 
    5719, 
    3175, 
    6533, 
    3494, 
    4328, 
    4525, 
    4101, 
    4048, 
    1477, 
    6531, 
    4349, 
    5747, 
    4048, 
    2404, 
    1477, 
    4272, 
    4048, 
    4101, 
    4164, 
    1893, 
    2404, 
    3916, 
    4164, 
    4048, 
    4894, 
    4328, 
    4117, 
    3916, 
    4718, 
    4164, 
    3916, 
    3646, 
    5275, 
    5275, 
    4525, 
    4718, 
    3916, 
    5275, 
    4718, 
    5747, 
    4349, 
    5275, 
    3646, 
    5747, 
    5275, 
    3646, 
    3341, 
    5747, 
    4164, 
    2404, 
    4048, 
    5234, 
    989, 
    1771, 
    4617, 
    4724, 
    5112, 
    4418, 
    4617, 
    2570, 
    4418, 
    4812, 
    4617, 
    2106, 
    989, 
    4548, 
    5020, 
    2764, 
    3609, 
    3175, 
    3494, 
    6533, 
    5675, 
    3005, 
    2764, 
    4349, 
    6531, 
    4137, 
    3341, 
    3005, 
    5675, 
    1488, 
    3851, 
    2106, 
    3090, 
    5956, 
    3131, 
    3134, 
    3090, 
    2715, 
    2772, 
    3417, 
    3090, 
    4349, 
    6533, 
    5275, 
    3778, 
    4328, 
    3494, 
    4894, 
    1158, 
    1893, 
    4328, 
    4894, 
    4718, 
    4117, 
    1158, 
    4894, 
    5020, 
    2823, 
    5719, 
    5886, 
    4965, 
    5650, 
    3609, 
    5886, 
    5650, 
    3303, 
    5106, 
    5886, 
    4418, 
    4206, 
    4812, 
    3306, 
    4206, 
    2965, 
    3306, 
    3978, 
    4206, 
    4240, 
    3175, 
    5642, 
    4011, 
    4240, 
    3712, 
    3494, 
    3175, 
    4240, 
    3778, 
    3494, 
    4011, 
    3134, 
    4039, 
    2772, 
    4164, 
    4894, 
    1893, 
    4039, 
    4117, 
    3778, 
    4039, 
    2203, 
    4117, 
    4718, 
    4894, 
    4164, 
    4328, 
    3778, 
    4117, 
    3303, 
    3741, 
    2962, 
    3134, 
    2715, 
    815, 
    5956, 
    2768, 
    3131, 
    3417, 
    5956, 
    3090, 
    3417, 
    2768, 
    5956, 
    4011, 
    3417, 
    2772, 
    3778, 
    4011, 
    2772, 
    3494, 
    4240, 
    4011, 
    3978, 
    5642, 
    4206, 
    3712, 
    3978, 
    3612, 
    3712, 
    4240, 
    5642, 
    3128, 
    3609, 
    2764, 
    2768, 
    6185, 
    3038, 
    3978, 
    3306, 
    3612, 
    2965, 
    2570, 
    4447, 
    4418, 
    2570, 
    2965, 
    2823, 
    4812, 
    4206, 
    4965, 
    5886, 
    5106, 
    4812, 
    4965, 
    4617, 
    5886, 
    3609, 
    3303, 
    4812, 
    5650, 
    4965, 
    4812, 
    5020, 
    5650, 
    2570, 
    4008, 
    4236, 
    2653, 
    2432, 
    2852, 
    759, 
    1595, 
    1901, 
    3851, 
    1855, 
    4457, 
    5444, 
    3851, 
    1488, 
    1108, 
    1855, 
    3851, 
    2577, 
    2051, 
    893, 
    3953, 
    2674, 
    3902, 
    4899, 
    3953, 
    3684, 
    2774, 
    5044, 
    3684, 
    3311, 
    3618, 
    4899, 
    4725, 
    1595, 
    2674, 
    4899, 
    4725, 
    3953, 
    3618, 
    2175, 
    4725, 
    4550, 
    2051, 
    2577, 
    2246, 
    1159, 
    2204, 
    2246, 
    1693, 
    1159, 
    3980, 
    4420, 
    2982, 
    3627, 
    1855, 
    1108, 
    5717, 
    3786, 
    1429, 
    2374, 
    5717, 
    1429, 
    4619, 
    3786, 
    5717, 
    2589, 
    4619, 
    3092, 
    4420, 
    5361, 
    4619, 
    2374, 
    1855, 
    3092, 
    4619, 
    5717, 
    2374, 
    2589, 
    4420, 
    4619, 
    3189, 
    2839, 
    3786, 
    1429, 
    2713, 
    5910, 
    893, 
    1894, 
    1693, 
    2190, 
    2564, 
    4214, 
    3941, 
    3671, 
    3515, 
    1335, 
    3941, 
    2321, 
    3455, 
    3671, 
    3941, 
    4179, 
    3866, 
    1716, 
    1254, 
    6041, 
    2264, 
    1317, 
    3866, 
    4179, 
    3866, 
    1317, 
    2307, 
    4739, 
    3866, 
    2307, 
    925, 
    1716, 
    3866, 
    1317, 
    4179, 
    1999, 
    4179, 
    1716, 
    2264, 
    2554, 
    2953, 
    689, 
    1716, 
    3596, 
    2526, 
    3596, 
    2070, 
    2839, 
    2710, 
    4445, 
    1608, 
    3625, 
    2658, 
    3042, 
    3221, 
    3625, 
    2871, 
    3319, 
    2658, 
    3625, 
    1318, 
    3319, 
    3221, 
    2000, 
    791, 
    5351, 
    4445, 
    773, 
    1608, 
    4234, 
    4445, 
    2710, 
    6256, 
    4359, 
    4675, 
    4234, 
    6256, 
    4445, 
    4234, 
    2453, 
    6256, 
    3894, 
    4146, 
    2453, 
    3674, 
    3944, 
    4359, 
    4532, 
    791, 
    1621, 
    3032, 
    4332, 
    2645, 
    4332, 
    5351, 
    4532, 
    5936, 
    3439, 
    2000, 
    5150, 
    5936, 
    1318, 
    5150, 
    2256, 
    5936, 
    4440, 
    1621, 
    2191, 
    3053, 
    4440, 
    2191, 
    2645, 
    4332, 
    4532, 
    1304, 
    2957, 
    1989, 
    4675, 
    4445, 
    6256, 
    4500, 
    4675, 
    4359, 
    1989, 
    773, 
    4675, 
    4480, 
    2295, 
    1759, 
    2980, 
    1939, 
    2957, 
    4480, 
    2980, 
    2295, 
    1229, 
    1939, 
    2980, 
    2957, 
    688, 
    5326, 
    2980, 
    2957, 
    1304, 
    1939, 
    688, 
    2957, 
    2295, 
    2980, 
    1304, 
    1229, 
    4848, 
    1939, 
    3091, 
    2746, 
    3113, 
    3248, 
    3558, 
    2716, 
    6117, 
    2751, 
    5096, 
    3979, 
    6117, 
    4207, 
    3979, 
    6004, 
    6117, 
    2651, 
    3979, 
    3037, 
    3713, 
    6004, 
    3979, 
    3831, 
    3444, 
    4097, 
    4097, 
    3444, 
    3117, 
    3091, 
    3831, 
    3418, 
    3091, 
    3558, 
    3831, 
    5451, 
    3762, 
    4027, 
    5451, 
    2778, 
    3762, 
    5375, 
    5451, 
    4027, 
    3444, 
    2778, 
    5451, 
    5451, 
    3117, 
    3444, 
    4253, 
    5375, 
    4027, 
    4253, 
    5278, 
    5375, 
    956, 
    1660, 
    1742, 
    2229, 
    1203, 
    970, 
    4598, 
    2229, 
    970, 
    2628, 
    2465, 
    2882, 
    4038, 
    1671, 
    2628, 
    1671, 
    861, 
    2628, 
    2819, 
    3924, 
    1412, 
    4038, 
    2628, 
    3015, 
    5795, 
    4038, 
    3015, 
    3775, 
    2229, 
    4038, 
    1909, 
    1877, 
    2366, 
    1188, 
    1909, 
    1845, 
    1877, 
    4300, 
    2366, 
    2060, 
    911, 
    5105, 
    2027, 
    747, 
    1974, 
    2284, 
    2027, 
    1287, 
    2907, 
    2284, 
    1287, 
    1979, 
    2951, 
    1287, 
    2492, 
    3315, 
    2907, 
    1287, 
    2951, 
    2907, 
    3072, 
    4854, 
    5008, 
    1460, 
    4369, 
    2392, 
    4632, 
    4809, 
    3017, 
    4367, 
    2527, 
    4564, 
    3907, 
    3583, 
    3277, 
    3262, 
    3907, 
    2920, 
    2581, 
    3583, 
    3907, 
    4709, 
    3273, 
    2931, 
    3277, 
    4709, 
    2935, 
    3277, 
    4541, 
    4709, 
    4291, 
    2828, 
    4072, 
    3579, 
    4291, 
    4072, 
    3595, 
    3291, 
    4498, 
    2692, 
    3595, 
    3579, 
    6486, 
    5872, 
    3909, 
    5997, 
    6486, 
    4158, 
    5997, 
    4575, 
    6486, 
    3595, 
    4498, 
    4291, 
    3291, 
    2951, 
    4674, 
    2907, 
    3291, 
    2492, 
    3333, 
    3639, 
    5778, 
    4884, 
    2527, 
    2935, 
    4709, 
    4884, 
    2935, 
    2931, 
    2522, 
    4884, 
    4884, 
    2522, 
    5153, 
    4709, 
    2931, 
    4884, 
    3579, 
    3273, 
    4541, 
    2492, 
    3595, 
    2692, 
    3595, 
    4291, 
    3579, 
    4072, 
    3179, 
    3809, 
    4072, 
    2828, 
    3179, 
    3273, 
    4072, 
    3809, 
    3273, 
    3579, 
    4072, 
    2492, 
    3291, 
    3595, 
    6160, 
    6441, 
    5499, 
    4156, 
    2508, 
    2920, 
    3907, 
    4156, 
    2920, 
    3277, 
    2935, 
    4156, 
    4618, 
    4883, 
    5035, 
    3418, 
    3713, 
    5433, 
    6109, 
    4463, 
    4644, 
    2542, 
    4463, 
    4253, 
    3178, 
    5857, 
    2996, 
    4644, 
    5089, 
    4820, 
    4947, 
    4041, 
    5089, 
    3979, 
    2651, 
    3713, 
    4207, 
    3037, 
    3979, 
    4207, 
    3369, 
    3037, 
    5278, 
    4463, 
    6109, 
    3117, 
    5375, 
    2751, 
    4253, 
    4463, 
    5278, 
    2451, 
    3369, 
    5035, 
    6109, 
    5096, 
    5278, 
    5046, 
    6109, 
    4644, 
    5046, 
    5367, 
    6109, 
    4707, 
    2522, 
    3532, 
    2869, 
    4707, 
    3219, 
    5153, 
    4728, 
    2527, 
    4883, 
    4787, 
    4707, 
    4618, 
    5269, 
    5171, 
    5096, 
    2751, 
    5278, 
    5269, 
    5367, 
    5046, 
    4207, 
    6117, 
    5096, 
    4787, 
    5153, 
    4707, 
    4657, 
    3265, 
    2923, 
    2451, 
    4477, 
    6344, 
    2451, 
    4268, 
    4477, 
    6344, 
    4477, 
    4657, 
    5742, 
    6344, 
    4657, 
    3369, 
    2451, 
    6344, 
    4475, 
    3387, 
    5343, 
    3287, 
    4656, 
    2947, 
    3683, 
    3387, 
    4475, 
    4656, 
    3683, 
    4475, 
    3593, 
    1892, 
    4832, 
    2403, 
    1474, 
    3952, 
    4504, 
    4686, 
    2098, 
    4686, 
    3683, 
    3952, 
    4685, 
    4505, 
    4504, 
    3194, 
    4685, 
    4504, 
    2844, 
    4853, 
    4685, 
    4301, 
    3387, 
    4505, 
    4207, 
    4419, 
    3369, 
    1742, 
    846, 
    2284, 
    846, 
    747, 
    2027, 
    61, 
    593, 
    4337, 
    593, 
    60, 
    1481, 
    4417, 
    4635, 
    723, 
    1509, 
    2614, 
    929, 
    1509, 
    2150, 
    2614, 
    1257, 
    1826, 
    856, 
    3300, 
    2391, 
    1444, 
    2639, 
    3300, 
    2959, 
    1876, 
    2391, 
    3300, 
    2959, 
    1444, 
    2080, 
    4172, 
    2959, 
    2080, 
    2639, 
    3025, 
    3300, 
    31, 
    6588, 
    1444, 
    3726, 
    734, 
    1571, 
    1492, 
    3726, 
    835, 
    1492, 
    2213, 
    3726, 
    2213, 
    1178, 
    1965, 
    734, 
    2213, 
    1965, 
    1492, 
    3453, 
    2213, 
    5448, 
    2760, 
    4893, 
    5672, 
    5116, 
    5239, 
    2543, 
    6530, 
    5239, 
    5477, 
    5957, 
    6450, 
    6530, 
    5477, 
    5672, 
    5239, 
    6530, 
    5672, 
    2543, 
    4633, 
    6530, 
    4810, 
    4961, 
    5957, 
    4975, 
    2760, 
    5116, 
    6389, 
    4007, 
    2765, 
    5116, 
    5672, 
    6450, 
    5957, 
    4961, 
    6291, 
    6450, 
    5957, 
    5654, 
    5477, 
    4810, 
    5957, 
    4822, 
    5978, 
    4975, 
    1492, 
    4822, 
    3453, 
    5978, 
    2760, 
    4975, 
    993, 
    3125, 
    5978, 
    5476, 
    6207, 
    3126, 
    2765, 
    1178, 
    2213, 
    334, 
    333, 
    5223, 
    6598, 
    64, 
    63, 
    1303, 
    6598, 
    63, 
    65, 
    64, 
    6598, 
    6691, 
    66, 
    65, 
    2294, 
    6691, 
    65, 
    67, 
    66, 
    6691, 
    68, 
    6691, 
    2294, 
    1303, 
    2294, 
    6598, 
    3878, 
    62, 
    883, 
    3878, 
    1303, 
    62, 
    888, 
    3878, 
    883, 
    6362, 
    2961, 
    5181, 
    2565, 
    5839, 
    3878, 
    2565, 
    2961, 
    5839, 
    67, 
    6691, 
    68, 
    65, 
    6598, 
    2294, 
    63, 
    62, 
    1303, 
    3878, 
    888, 
    2565, 
    5331, 
    2407, 
    1895, 
    5231, 
    5331, 
    3325, 
    5231, 
    4537, 
    5331, 
    4337, 
    4537, 
    883, 
    4337, 
    593, 
    4537, 
    1935, 
    1220, 
    4381, 
    1827, 
    1935, 
    676, 
    3466, 
    1163, 
    2206, 
    4381, 
    3466, 
    2206, 
    1645, 
    4381, 
    2206, 
    3261, 
    1935, 
    4381, 
    1220, 
    2988, 
    3466, 
    2988, 
    3325, 
    3466, 
    2988, 
    5231, 
    3325, 
    4019, 
    1397, 
    3753, 
    3325, 
    5331, 
    1895, 
    1163, 
    3325, 
    1895, 
    5231, 
    888, 
    883, 
    1481, 
    5331, 
    4537, 
    2988, 
    888, 
    5231, 
    5107, 
    4966, 
    1481, 
    4019, 
    5107, 
    1397, 
    4019, 
    4249, 
    5107, 
    730, 
    1481, 
    60, 
    4249, 
    4966, 
    5107, 
    3753, 
    1262, 
    1830, 
    3753, 
    1397, 
    1262, 
    1075, 
    5177, 
    1830, 
    1481, 
    4966, 
    2407, 
    6419, 
    6123, 
    5521, 
    4019, 
    6419, 
    5521, 
    6228, 
    6123, 
    6419, 
    5177, 
    6228, 
    6400, 
    5177, 
    2576, 
    6228, 
    4966, 
    4456, 
    2407, 
    5521, 
    4249, 
    4019, 
    6400, 
    6228, 
    6419, 
    3753, 
    6400, 
    4019, 
    3753, 
    1830, 
    6400, 
    6219, 
    5333, 
    5236, 
    4249, 
    6219, 
    4456, 
    5850, 
    5333, 
    6219, 
    6123, 
    5850, 
    5521, 
    2572, 
    4722, 
    5850, 
    4456, 
    4640, 
    1895, 
    5850, 
    4722, 
    5333, 
    4897, 
    4327, 
    4523, 
    5333, 
    4722, 
    4897, 
    5236, 
    5333, 
    4897, 
    6219, 
    4249, 
    5521, 
    5557, 
    3846, 
    4113, 
    4722, 
    5557, 
    5220, 
    2572, 
    2967, 
    5557, 
    4942, 
    1382, 
    2346, 
    730, 
    4942, 
    1397, 
    730, 
    59, 
    4942, 
    59, 
    730, 
    60, 
    4792, 
    39, 
    592, 
    36, 
    4792, 
    37, 
    4818, 
    2576, 
    39, 
    4642, 
    4818, 
    4792, 
    4642, 
    5703, 
    4818, 
    5220, 
    4113, 
    4327, 
    4897, 
    5220, 
    4327, 
    4722, 
    2572, 
    5557, 
    4640, 
    5236, 
    1163, 
    5220, 
    4897, 
    4722, 
    5236, 
    2206, 
    1163, 
    4523, 
    4950, 
    4897, 
    4523, 
    1645, 
    4950, 
    4907, 
    5050, 
    3323, 
    1262, 
    869, 
    43, 
    1830, 
    1262, 
    43, 
    5557, 
    6192, 
    3846, 
    5874, 
    6228, 
    3457, 
    3745, 
    5874, 
    3457, 
    6400, 
    6419, 
    4019, 
    5733, 
    6123, 
    5874, 
    5733, 
    5850, 
    6123, 
    3307, 
    5961, 
    6192, 
    5874, 
    6123, 
    6228, 
    2967, 
    5733, 
    5663, 
    2572, 
    5850, 
    5733, 
    2770, 
    929, 
    3614, 
    5107, 
    730, 
    1397, 
    4456, 
    4966, 
    4249, 
    1481, 
    730, 
    5107, 
    1075, 
    2576, 
    5177, 
    4327, 
    2575, 
    2970, 
    5557, 
    4113, 
    5220, 
    4559, 
    3900, 
    4149, 
    6192, 
    2513, 
    3846, 
    2967, 
    6192, 
    5557, 
    2967, 
    3307, 
    6192, 
    4907, 
    3632, 
    4736, 
    5863, 
    4907, 
    4736, 
    3846, 
    5863, 
    4736, 
    3846, 
    2513, 
    5863, 
    6287, 
    2924, 
    5050, 
    4907, 
    6287, 
    5050, 
    2513, 
    2924, 
    6287, 
    1397, 
    869, 
    1262, 
    4212, 
    3613, 
    2623, 
    1223, 
    4262, 
    1937, 
    2815, 
    3613, 
    3883, 
    3169, 
    3010, 
    3613, 
    1086, 
    3010, 
    1838, 
    4985, 
    4746, 
    5244, 
    1086, 
    4985, 
    3010, 
    1086, 
    2159, 
    4985, 
    1537, 
    680, 
    4212, 
    4661, 
    1537, 
    4212, 
    5244, 
    4918, 
    4661, 
    4985, 
    5244, 
    2623, 
    4746, 
    4918, 
    5244, 
    2130, 
    1537, 
    4661, 
    4746, 
    3165, 
    3484, 
    3010, 
    4985, 
    2623, 
    2159, 
    3165, 
    4746, 
    1035, 
    4650, 
    4816, 
    4650, 
    1098, 
    1847, 
    4816, 
    4650, 
    1847, 
    2368, 
    4816, 
    1847, 
    2130, 
    1035, 
    4816, 
    1035, 
    1801, 
    4650, 
    6122, 
    6499, 
    3484, 
    6499, 
    2338, 
    1801, 
    1035, 
    3484, 
    6499, 
    2460, 
    2603, 
    2537, 
    1967, 
    2460, 
    736, 
    1967, 
    1266, 
    2993, 
    5354, 
    1584, 
    2169, 
    5325, 
    736, 
    2460, 
    2537, 
    5325, 
    2460, 
    3165, 
    1572, 
    5325, 
    1364, 
    4574, 
    2338, 
    3236, 
    1049, 
    1810, 
    6505, 
    3615, 
    3308, 
    2578, 
    5043, 
    2972, 
    3884, 
    3615, 
    4898, 
    1213, 
    3884, 
    5043, 
    1213, 
    1929, 
    3884, 
    2139, 
    1049, 
    2459, 
    4208, 
    2139, 
    2459, 
    1547, 
    2368, 
    2139, 
    1416, 
    1547, 
    694, 
    2368, 
    1847, 
    2139, 
    1416, 
    2368, 
    1547, 
    4120, 
    1537, 
    2130, 
    1416, 
    4120, 
    2368, 
    1416, 
    4426, 
    4120, 
    5354, 
    2338, 
    4574, 
    1098, 
    5500, 
    2169, 
    1801, 
    2338, 
    5354, 
    2681, 
    1384, 
    2038, 
    872, 
    2876, 
    2038, 
    5261, 
    5154, 
    2505, 
    2876, 
    3061, 
    2681, 
    5261, 
    2505, 
    2917, 
    3076, 
    5154, 
    2700, 
    3076, 
    5017, 
    5154, 
    3061, 
    5805, 
    2700, 
    4867, 
    3703, 
    4694, 
    1098, 
    1810, 
    1049, 
    4106, 
    3196, 
    2847, 
    3792, 
    3512, 
    3567, 
    2036, 
    3792, 
    3567, 
    862, 
    1672, 
    5349, 
    2648, 
    2644, 
    3512, 
    4943, 
    1384, 
    2681, 
    4104, 
    1810, 
    2344, 
    2459, 
    3236, 
    2892, 
    2459, 
    1049, 
    3236, 
    2169, 
    2344, 
    1810, 
    1584, 
    1374, 
    2344, 
    1847, 
    1098, 
    1049, 
    4120, 
    2130, 
    4816, 
    2368, 
    4120, 
    4816, 
    3757, 
    819, 
    2014, 
    2985, 
    3757, 
    2014, 
    1534, 
    676, 
    3757, 
    5950, 
    3801, 
    4971, 
    3884, 
    1929, 
    2439, 
    1213, 
    1881, 
    1929, 
    5161, 
    2718, 
    3888, 
    4404, 
    2459, 
    2892, 
    2476, 
    4404, 
    2892, 
    4190, 
    4292, 
    4404, 
    872, 
    959, 
    2094, 
    1681, 
    872, 
    2094, 
    5263, 
    4292, 
    5161, 
    2529, 
    5770, 
    4190, 
    5770, 
    3814, 
    4076, 
    4190, 
    5770, 
    4076, 
    2529, 
    3690, 
    5770, 
    2139, 
    1847, 
    1049, 
    1945, 
    2063, 
    694, 
    4426, 
    1537, 
    4120, 
    750, 
    1977, 
    2036, 
    5370, 
    4624, 
    5319, 
    872, 
    2038, 
    959, 
    2504, 
    2006, 
    805, 
    1384, 
    2287, 
    1745, 
    2927, 
    1329, 
    2006, 
    2504, 
    2927, 
    2006, 
    6055, 
    2516, 
    1981, 
    4302, 
    6055, 
    4087, 
    4423, 
    2516, 
    6055, 
    2916, 
    3268, 
    2927, 
    2916, 
    3258, 
    3268, 
    4423, 
    3268, 
    2516, 
    2315, 
    4423, 
    4302, 
    2927, 
    3268, 
    4423, 
    1290, 
    1981, 
    2516, 
    4677, 
    5158, 
    3659, 
    5139, 
    3470, 
    1856, 
    5158, 
    3357, 
    3659, 
    6036, 
    5158, 
    4677, 
    1908, 
    3357, 
    5158, 
    3470, 
    2375, 
    1856, 
    3827, 
    1430, 
    2375, 
    3470, 
    3827, 
    2375, 
    1243, 
    2257, 
    3827, 
    2807, 
    896, 
    2562, 
    6213, 
    2053, 
    1403, 
    1469, 
    896, 
    2053, 
    3492, 
    2821, 
    4747, 
    3651, 
    3776, 
    3347, 
    2450, 
    4198, 
    3347, 
    3921, 
    969, 
    4858, 
    5149, 
    2821, 
    3492, 
    5012, 
    5149, 
    3492, 
    2680, 
    3060, 
    5149, 
    3486, 
    3770, 
    3167, 
    2813, 
    2868, 
    2394, 
    1403, 
    969, 
    6213, 
    2868, 
    1881, 
    2394, 
    3012, 
    2868, 
    2450, 
    1144, 
    1881, 
    2868, 
    1144, 
    1929, 
    1881, 
    1929, 
    1144, 
    665, 
    4798, 
    1463, 
    2094, 
    3793, 
    2813, 
    1463, 
    959, 
    4798, 
    2094, 
    3167, 
    2813, 
    3793, 
    1888, 
    3486, 
    4624, 
    3966, 
    2398, 
    1469, 
    3167, 
    3770, 
    5937, 
    3486, 
    1888, 
    3770, 
    4433, 
    3486, 
    3167, 
    1888, 
    2398, 
    3770, 
    2450, 
    2868, 
    2813, 
    1213, 
    2394, 
    1881, 
    1213, 
    2235, 
    2394, 
    3856, 
    2348, 
    5221, 
    1384, 
    3856, 
    2287, 
    1384, 
    2348, 
    3856, 
    1888, 
    1152, 
    2248, 
    2813, 
    2394, 
    1463, 
    2450, 
    2813, 
    3167, 
    3258, 
    2287, 
    1290, 
    3447, 
    3258, 
    2916, 
    5700, 
    3447, 
    2916, 
    2504, 
    5700, 
    2916, 
    2754, 
    3447, 
    5700, 
    3121, 
    1745, 
    3447, 
    1745, 
    2287, 
    3258, 
    4726, 
    4103, 
    1944, 
    5045, 
    4516, 
    4726, 
    2896, 
    5085, 
    2480, 
    4353, 
    4516, 
    5045, 
    4353, 
    3837, 
    4516, 
    2198, 
    1944, 
    1234, 
    1632, 
    693, 
    1944, 
    2315, 
    1047, 
    1329, 
    2315, 
    1778, 
    1808, 
    2927, 
    4423, 
    1329, 
    4087, 
    760, 
    2586, 
    3495, 
    3939, 
    2034, 
    1778, 
    2342, 
    1808, 
    1001, 
    1372, 
    2342, 
    5372, 
    2586, 
    2176, 
    1109, 
    5372, 
    2176, 
    5272, 
    2979, 
    5372, 
    1001, 
    2979, 
    5272, 
    5139, 
    1551, 
    708, 
    1596, 
    4224, 
    2176, 
    1596, 
    4627, 
    4224, 
    4627, 
    2143, 
    4224, 
    760, 
    4627, 
    1596, 
    4506, 
    2143, 
    4627, 
    4224, 
    1109, 
    2176, 
    6030, 
    3495, 
    860, 
    2749, 
    4637, 
    2555, 
    5932, 
    3495, 
    6030, 
    4637, 
    5932, 
    4452, 
    3176, 
    3495, 
    5932, 
    5288, 
    3301, 
    2108, 
    1494, 
    5288, 
    2108, 
    2807, 
    2562, 
    5288, 
    2398, 
    1888, 
    1697, 
    1469, 
    2398, 
    896, 
    4198, 
    3651, 
    3347, 
    5937, 
    4198, 
    2450, 
    3167, 
    5937, 
    2450, 
    3770, 
    3966, 
    5937, 
    6111, 
    3651, 
    4198, 
    3966, 
    6111, 
    4198, 
    3966, 
    6213, 
    6111, 
    2398, 
    3966, 
    3770, 
    6213, 
    3921, 
    6111, 
    1469, 
    6213, 
    3966, 
    1469, 
    2053, 
    6213, 
    3301, 
    1774, 
    996, 
    2108, 
    3301, 
    996, 
    2562, 
    1697, 
    3607, 
    2198, 
    1234, 
    1152, 
    4624, 
    4433, 
    5319, 
    1888, 
    4624, 
    1152, 
    3486, 
    4433, 
    4624, 
    1632, 
    1944, 
    2198, 
    4798, 
    959, 
    3121, 
    805, 
    693, 
    1632, 
    2510, 
    798, 
    2788, 
    5085, 
    5045, 
    2480, 
    2004, 
    5085, 
    2896, 
    4353, 
    5045, 
    5085, 
    2312, 
    4353, 
    1324, 
    3837, 
    4103, 
    4516, 
    5313, 
    1545, 
    3518, 
    5045, 
    5313, 
    2480, 
    4726, 
    693, 
    5313, 
    5349, 
    5630, 
    2648, 
    3792, 
    5349, 
    2648, 
    6446, 
    1736, 
    5793, 
    5139, 
    4224, 
    1551, 
    3470, 
    5139, 
    708, 
    1109, 
    4224, 
    5139, 
    4052, 
    1059, 
    3259, 
    4224, 
    2143, 
    1551, 
    4694, 
    4106, 
    2705, 
    2476, 
    4517, 
    3703, 
    4201, 
    4321, 
    5471, 
    3236, 
    4201, 
    2892, 
    4104, 
    4107, 
    4321, 
    5394, 
    2709, 
    3085, 
    2644, 
    5512, 
    3031, 
    2485, 
    2709, 
    5297, 
    3690, 
    5749, 
    3393, 
    2476, 
    3703, 
    2529, 
    5154, 
    5413, 
    2505, 
    2847, 
    3031, 
    3363, 
    4106, 
    2847, 
    2705, 
    3841, 
    3567, 
    3512, 
    4106, 
    3841, 
    3196, 
    4694, 
    4517, 
    5471, 
    3081, 
    4867, 
    5935, 
    3703, 
    4517, 
    4694, 
    4517, 
    2476, 
    2892, 
    4201, 
    3236, 
    4104, 
    3512, 
    2644, 
    3196, 
    5394, 
    5297, 
    2709, 
    3412, 
    5466, 
    3085, 
    6351, 
    6076, 
    5394, 
    3196, 
    3031, 
    2847, 
    5512, 
    2485, 
    5297, 
    6076, 
    5512, 
    5297, 
    5394, 
    6076, 
    5297, 
    3363, 
    3031, 
    6076, 
    2644, 
    5843, 
    6418, 
    5359, 
    5261, 
    2917, 
    2348, 
    5359, 
    1816, 
    4943, 
    5261, 
    5359, 
    4586, 
    4387, 
    4175, 
    3789, 
    4758, 
    3508, 
    4052, 
    3972, 
    4586, 
    2505, 
    3707, 
    2917, 
    5298, 
    3664, 
    3935, 
    4943, 
    5359, 
    2348, 
    1551, 
    4758, 
    3789, 
    2917, 
    3972, 
    3259, 
    4387, 
    3935, 
    4175, 
    1059, 
    1816, 
    3259, 
    2518, 
    331, 
    632, 
    2929, 
    875, 
    2040, 
    1387, 
    3437, 
    2040, 
    1965, 
    5223, 
    2929, 
    3726, 
    2213, 
    734, 
    1178, 
    5223, 
    1965, 
    332, 
    331, 
    875, 
    4337, 
    62, 
    61, 
    1481, 
    4537, 
    593, 
    883, 
    62, 
    4337, 
    1481, 
    2407, 
    5331, 
    6285, 
    1827, 
    5525, 
    3950, 
    1276, 
    2279, 
    2961, 
    3950, 
    2279, 
    2565, 
    2048, 
    4396, 
    883, 
    4537, 
    5231, 
    5339, 
    5525, 
    6515, 
    4396, 
    5339, 
    6515, 
    1220, 
    1935, 
    6285, 
    6362, 
    5839, 
    2961, 
    2294, 
    6362, 
    5181, 
    2294, 
    1303, 
    6362, 
    1793, 
    685, 
    136, 
    4121, 
    1538, 
    683, 
    1585, 
    4121, 
    683, 
    751, 
    1538, 
    4121, 
    927, 
    685, 
    1538, 
    3926, 
    2631, 
    5916, 
    3926, 
    2794, 
    2631, 
    1279, 
    3926, 
    2786, 
    3151, 
    2794, 
    3926, 
    1585, 
    4562, 
    751, 
    4562, 
    4830, 
    5191, 
    4264, 
    5052, 
    2794, 
    1279, 
    685, 
    927, 
    2518, 
    2040, 
    875, 
    1562, 
    2490, 
    722, 
    6172, 
    2040, 
    2518, 
    3378, 
    2149, 
    1562, 
    722, 
    5184, 
    1562, 
    3045, 
    2661, 
    5597, 
    5184, 
    3045, 
    3378, 
    1562, 
    5184, 
    3378, 
    722, 
    330, 
    5314, 
    5597, 
    5423, 
    2601, 
    3904, 
    5597, 
    3636, 
    2661, 
    5423, 
    5597, 
    327, 
    2661, 
    631, 
    5744, 
    2991, 
    3329, 
    5314, 
    329, 
    328, 
    2663, 
    1236, 
    2251, 
    5744, 
    3636, 
    5597, 
    2991, 
    5744, 
    2601, 
    3329, 
    3636, 
    5744, 
    696, 
    3329, 
    2991, 
    4594, 
    3379, 
    4394, 
    696, 
    1484, 
    4421, 
    5423, 
    325, 
    2601, 
    902, 
    2991, 
    4365, 
    4365, 
    325, 
    324, 
    4766, 
    2663, 
    4594, 
    5423, 
    326, 
    325, 
    5744, 
    5597, 
    2601, 
    327, 
    326, 
    5423, 
    4154, 
    3378, 
    5855, 
    5053, 
    4154, 
    3904, 
    6176, 
    5053, 
    3904, 
    4184, 
    1071, 
    5053, 
    2149, 
    3378, 
    4154, 
    4577, 
    324, 
    323, 
    1484, 
    696, 
    902, 
    6288, 
    2820, 
    4043, 
    2251, 
    3173, 
    6288, 
    2251, 
    1236, 
    3173, 
    2691, 
    5488, 
    985, 
    2104, 
    2691, 
    985, 
    3781, 
    3491, 
    2022, 
    4266, 
    4311, 
    2902, 
    4410, 
    1655, 
    840, 
    5766, 
    3044, 
    2487, 
    6047, 
    5766, 
    2902, 
    3377, 
    3044, 
    5766, 
    6047, 
    3676, 
    3377, 
    3491, 
    3781, 
    3243, 
    2022, 
    1358, 
    3781, 
    4138, 
    5145, 
    1795, 
    6047, 
    3781, 
    3676, 
    5766, 
    6047, 
    3377, 
    3243, 
    3781, 
    6047, 
    1358, 
    2334, 
    3676, 
    4836, 
    3305, 
    1617, 
    2660, 
    4836, 
    786, 
    2660, 
    3044, 
    5126, 
    3305, 
    2964, 
    2187, 
    5419, 
    4587, 
    2569, 
    4138, 
    5233, 
    3881, 
    2125, 
    1531, 
    4759, 
    4932, 
    1531, 
    3974, 
    2942, 
    865, 
    1455, 
    5966, 
    3283, 
    2942, 
    4879, 
    5966, 
    2942, 
    4879, 
    5029, 
    5966, 
    4308, 
    4879, 
    2684, 
    4092, 
    3826, 
    5029, 
    3918, 
    2769, 
    3197, 
    5763, 
    3918, 
    3197, 
    2848, 
    5812, 
    3197, 
    3386, 
    3529, 
    5763, 
    6065, 
    3217, 
    4186, 
    5763, 
    6065, 
    3918, 
    3529, 
    3217, 
    6065, 
    4398, 
    3456, 
    5776, 
    2866, 
    4398, 
    4186, 
    1086, 
    1838, 
    4398, 
    3386, 
    6359, 
    2942, 
    5276, 
    3152, 
    1617, 
    2769, 
    5176, 
    3197, 
    2796, 
    3152, 
    5176, 
    6359, 
    1873, 
    865, 
    2848, 
    6359, 
    5812, 
    1134, 
    1873, 
    6359, 
    2964, 
    1134, 
    2187, 
    1617, 
    3305, 
    2187, 
    4388, 
    2802, 
    1873, 
    2569, 
    4388, 
    2964, 
    5397, 
    4932, 
    3974, 
    2802, 
    5397, 
    3157, 
    4587, 
    4932, 
    5397, 
    2569, 
    4587, 
    4388, 
    5419, 
    3881, 
    5233, 
    1966, 
    2125, 
    1028, 
    3974, 
    672, 
    3477, 
    735, 
    1531, 
    2125, 
    5397, 
    3974, 
    3157, 
    4759, 
    4932, 
    4587, 
    4759, 
    1531, 
    4932, 
    4879, 
    2942, 
    1455, 
    3861, 
    3529, 
    3590, 
    3529, 
    6065, 
    5763, 
    4186, 
    4165, 
    6065, 
    2448, 
    4398, 
    2866, 
    5776, 
    3132, 
    4165, 
    4398, 
    5776, 
    4186, 
    3456, 
    3132, 
    5776, 
    6359, 
    2848, 
    1134, 
    3386, 
    5812, 
    6359, 
    3386, 
    5763, 
    5812, 
    3529, 
    3386, 
    3283, 
    3590, 
    3529, 
    3283, 
    5966, 
    5029, 
    5711, 
    5364, 
    3240, 
    2900, 
    5266, 
    5364, 
    4125, 
    5266, 
    3240, 
    5364, 
    4165, 
    3132, 
    2769, 
    6065, 
    4165, 
    3918, 
    3217, 
    2866, 
    4186, 
    5763, 
    3197, 
    5812, 
    6077, 
    5176, 
    2769, 
    4948, 
    6077, 
    2769, 
    2796, 
    5176, 
    6077, 
    3386, 
    2942, 
    3283, 
    1937, 
    4262, 
    3883, 
    5416, 
    1825, 
    2354, 
    2763, 
    886, 
    1691, 
    3127, 
    2763, 
    5274, 
    711, 
    3127, 
    1952, 
    711, 
    1553, 
    4710, 
    2047, 
    886, 
    2763, 
    5076, 
    2047, 
    2763, 
    5469, 
    5076, 
    3127, 
    711, 
    5469, 
    3127, 
    4710, 
    4542, 
    5469, 
    4542, 
    1395, 
    5076, 
    4184, 
    2354, 
    1825, 
    4184, 
    3948, 
    2354, 
    1071, 
    4184, 
    1825, 
    5053, 
    4394, 
    4184, 
    3677, 
    3601, 
    3948, 
    2517, 
    3870, 
    3379, 
    3601, 
    1395, 
    3948, 
    2145, 
    2547, 
    1553, 
    5855, 
    3904, 
    4154, 
    5597, 
    5855, 
    3045, 
    5597, 
    3904, 
    5855, 
    6273, 
    4594, 
    6176, 
    1946, 
    4766, 
    3329, 
    1946, 
    1236, 
    4766, 
    3379, 
    3677, 
    4394, 
    2663, 
    2251, 
    2928, 
    3181, 
    3500, 
    2493, 
    4184, 
    3677, 
    3948, 
    2820, 
    1766, 
    698, 
    4269, 
    4043, 
    2820, 
    1313, 
    4269, 
    698, 
    1313, 
    1996, 
    4478, 
    4421, 
    1236, 
    1946, 
    1766, 
    3247, 
    985, 
    3173, 
    1236, 
    3247, 
    2928, 
    2251, 
    1700, 
    900, 
    4348, 
    1700, 
    2517, 
    3379, 
    2928, 
    900, 
    3500, 
    4348, 
    2047, 
    1395, 
    3601, 
    3173, 
    3247, 
    2820, 
    3783, 
    4043, 
    5124, 
    2241, 
    1223, 
    3488, 
    2831, 
    3559, 
    1691, 
    3169, 
    1406, 
    2360, 
    2063, 
    1416, 
    694, 
    914, 
    2063, 
    1945, 
    914, 
    5209, 
    2063, 
    2250, 
    1708, 
    1235, 
    4139, 
    4817, 
    1235, 
    1945, 
    4139, 
    1235, 
    1929, 
    665, 
    2439, 
    1698, 
    2259, 
    2250, 
    1952, 
    1245, 
    898, 
    2055, 
    1952, 
    898, 
    3127, 
    5076, 
    2763, 
    2259, 
    3832, 
    3488, 
    2763, 
    1691, 
    3832, 
    5222, 
    4547, 
    4717, 
    4426, 
    1416, 
    2063, 
    5209, 
    4426, 
    2063, 
    680, 
    1537, 
    4426, 
    4348, 
    2517, 
    2928, 
    1700, 
    4348, 
    2928, 
    3500, 
    3181, 
    4547, 
    2056, 
    3500, 
    900, 
    3500, 
    4547, 
    4348, 
    3249, 
    3181, 
    2493, 
    3772, 
    3249, 
    2493, 
    4262, 
    1223, 
    2241, 
    3249, 
    6336, 
    3559, 
    2815, 
    3883, 
    4262, 
    5222, 
    886, 
    2047, 
    3601, 
    5222, 
    2047, 
    4547, 
    3181, 
    4717, 
    2104, 
    985, 
    3247, 
    1484, 
    2104, 
    4421, 
    4096, 
    686, 
    1539, 
    4096, 
    3295, 
    686, 
    2133, 
    5260, 
    1539, 
    5922, 
    3963, 
    4513, 
    4513, 
    3602, 
    4313, 
    2104, 
    3871, 
    2691, 
    2104, 
    1484, 
    3871, 
    1484, 
    902, 
    5063, 
    4577, 
    902, 
    324, 
    4926, 
    4577, 
    323, 
    1228, 
    4926, 
    323, 
    3295, 
    3602, 
    4926, 
    4926, 
    5063, 
    4577, 
    3247, 
    1766, 
    2820, 
    3492, 
    3776, 
    5012, 
    6154, 
    1603, 
    4546, 
    5476, 
    2761, 
    4893, 
    993, 
    6207, 
    3125, 
    3126, 
    2761, 
    5476, 
    6207, 
    1353, 
    2310, 
    3125, 
    6207, 
    5476, 
    993, 
    1353, 
    6207, 
    2310, 
    1321, 
    3126, 
    3876, 
    3608, 
    5745, 
    1321, 
    5230, 
    3126, 
    5230, 
    2002, 
    4346, 
    4346, 
    3060, 
    2680, 
    5230, 
    4346, 
    5560, 
    3126, 
    5230, 
    3876, 
    1321, 
    2002, 
    5230, 
    2002, 
    3060, 
    4346, 
    1298, 
    1570, 
    5574, 
    5476, 
    2760, 
    3125, 
    5560, 
    4346, 
    2680, 
    4716, 
    5560, 
    2680, 
    3608, 
    3876, 
    5560, 
    6034, 
    6154, 
    5745, 
    4430, 
    1603, 
    732, 
    5407, 
    4430, 
    732, 
    1355, 
    1603, 
    4430, 
    6161, 
    5448, 
    4893, 
    4546, 
    6324, 
    4715, 
    5239, 
    5448, 
    6161, 
    2543, 
    5239, 
    5273, 
    2021, 
    1355, 
    4430, 
    5407, 
    2021, 
    4430, 
    1570, 
    5407, 
    732, 
    1570, 
    5040, 
    5407, 
    837, 
    2845, 
    4823, 
    4823, 
    2021, 
    837, 
    4976, 
    3946, 
    4823, 
    3390, 
    4182, 
    1579, 
    6083, 
    3057, 
    1355, 
    3390, 
    6083, 
    4182, 
    3390, 
    3057, 
    6083, 
    6083, 
    1355, 
    3946, 
    1603, 
    1355, 
    1263, 
    4182, 
    745, 
    1579, 
    1025, 
    933, 
    1863, 
    2464, 
    3726, 
    1571, 
    4975, 
    6084, 
    4822, 
    336, 
    4007, 
    2243, 
    6389, 
    3453, 
    4822, 
    6207, 
    2310, 
    3126, 
    5273, 
    1263, 
    1117, 
    2500, 
    1571, 
    3437, 
    1818, 
    2500, 
    2350, 
    2157, 
    1571, 
    2500, 
    2464, 
    1571, 
    2157, 
    1084, 
    5291, 
    2157, 
    835, 
    3726, 
    2464, 
    734, 
    3437, 
    1571, 
    2055, 
    1405, 
    711, 
    3642, 
    2123, 
    1024, 
    3865, 
    3642, 
    1024, 
    6080, 
    3865, 
    1024, 
    2002, 
    6080, 
    1024, 
    2699, 
    3865, 
    6080, 
    2545, 
    4341, 
    3865, 
    3336, 
    4374, 
    4566, 
    4160, 
    4374, 
    3000, 
    4566, 
    1526, 
    2123, 
    898, 
    2612, 
    2055, 
    2002, 
    1024, 
    795, 
    5574, 
    2563, 
    1298, 
    5745, 
    6154, 
    5449, 
    3126, 
    3876, 
    2761, 
    5560, 
    4716, 
    3608, 
    4716, 
    2563, 
    3302, 
    3608, 
    4716, 
    3302, 
    5012, 
    3776, 
    4858, 
    5590, 
    5012, 
    4858, 
    2680, 
    5149, 
    5012, 
    1624, 
    2821, 
    795, 
    1624, 
    2194, 
    4747, 
    1321, 
    6080, 
    2002, 
    3876, 
    5230, 
    5560, 
    795, 
    3060, 
    2002, 
    795, 
    2821, 
    3060, 
    2437, 
    5291, 
    1837, 
    2699, 
    2310, 
    2857, 
    5291, 
    2464, 
    2157, 
    993, 
    3739, 
    5386, 
    993, 
    835, 
    3739, 
    3135, 
    3101, 
    1062, 
    2350, 
    5215, 
    1818, 
    2773, 
    3101, 
    3135, 
    1825, 
    2729, 
    1071, 
    2547, 
    2145, 
    3101, 
    3101, 
    2145, 
    1062, 
    5416, 
    2547, 
    2729, 
    1825, 
    5416, 
    2729, 
    2354, 
    4542, 
    5416, 
    2354, 
    1395, 
    4542, 
    2831, 
    886, 
    4717, 
    2354, 
    3948, 
    1395, 
    4547, 
    2517, 
    4348, 
    2831, 
    4717, 
    3181, 
    6167, 
    2517, 
    4547, 
    5222, 
    6167, 
    4547, 
    3870, 
    2517, 
    6167, 
    3677, 
    3870, 
    3601, 
    3677, 
    3379, 
    3870, 
    5053, 
    1071, 
    4154, 
    2663, 
    2928, 
    3379, 
    5855, 
    3378, 
    3045, 
    6176, 
    3904, 
    3636, 
    6176, 
    4394, 
    5053, 
    6273, 
    6176, 
    3636, 
    4594, 
    4394, 
    6176, 
    6273, 
    4766, 
    4594, 
    3329, 
    6273, 
    3636, 
    3329, 
    4766, 
    6273, 
    2663, 
    3379, 
    4594, 
    3677, 
    4184, 
    4394, 
    1071, 
    2149, 
    4154, 
    4766, 
    1236, 
    2663, 
    4710, 
    1553, 
    2547, 
    5416, 
    4710, 
    2547, 
    4542, 
    5076, 
    5469, 
    5416, 
    4542, 
    4710, 
    1395, 
    2047, 
    5076, 
    1553, 
    2359, 
    2145, 
    1405, 
    1553, 
    711, 
    1837, 
    1084, 
    5058, 
    2359, 
    1837, 
    2145, 
    1405, 
    2359, 
    1553, 
    2699, 
    6080, 
    1321, 
    2950, 
    2545, 
    5441, 
    5402, 
    2950, 
    5441, 
    1837, 
    5402, 
    2437, 
    1837, 
    2359, 
    5402, 
    2359, 
    1405, 
    3290, 
    4130, 
    3290, 
    1405, 
    3000, 
    4130, 
    2612, 
    3000, 
    3336, 
    4341, 
    2699, 
    2545, 
    3865, 
    2310, 
    2699, 
    1321, 
    2310, 
    1353, 
    2857, 
    5386, 
    1353, 
    993, 
    5386, 
    2857, 
    1353, 
    2464, 
    5386, 
    3739, 
    5291, 
    2857, 
    5386, 
    2464, 
    5291, 
    5386, 
    1084, 
    1837, 
    5291, 
    2437, 
    5441, 
    2857, 
    2359, 
    2950, 
    5402, 
    2612, 
    4130, 
    2055, 
    3739, 
    835, 
    2464, 
    2055, 
    711, 
    1952, 
    5441, 
    2699, 
    2857, 
    5402, 
    5441, 
    2437, 
    2545, 
    2699, 
    5441, 
    1837, 
    1062, 
    2145, 
    5058, 
    1062, 
    1837, 
    2157, 
    2500, 
    5058, 
    2437, 
    2857, 
    5291, 
    2500, 
    1387, 
    2350, 
    2793, 
    2490, 
    1562, 
    6187, 
    2793, 
    2149, 
    1071, 
    6187, 
    2149, 
    2773, 
    3135, 
    6187, 
    6187, 
    3135, 
    5215, 
    1965, 
    2929, 
    734, 
    2350, 
    1387, 
    3733, 
    5058, 
    2500, 
    1818, 
    1062, 
    5058, 
    1818, 
    1084, 
    2157, 
    5058, 
    3733, 
    2490, 
    2793, 
    5215, 
    3733, 
    2793, 
    6187, 
    5215, 
    2793, 
    3135, 
    1818, 
    5215, 
    1387, 
    2040, 
    6172, 
    2793, 
    1562, 
    2149, 
    4183, 
    328, 
    631, 
    3045, 
    4183, 
    2661, 
    3045, 
    5184, 
    4183, 
    711, 
    4710, 
    5469, 
    3101, 
    2773, 
    2729, 
    2547, 
    3101, 
    2729, 
    1062, 
    1818, 
    3135, 
    5423, 
    2661, 
    327, 
    2773, 
    6187, 
    1071, 
    2729, 
    2773, 
    1071, 
    5215, 
    2350, 
    3733, 
    4183, 
    5184, 
    5314, 
    5314, 
    5184, 
    722, 
    329, 
    5314, 
    330, 
    328, 
    4183, 
    5314, 
    4183, 
    631, 
    2661, 
    5209, 
    1937, 
    680, 
    3488, 
    5209, 
    914, 
    3488, 
    1223, 
    5209, 
    5209, 
    1223, 
    1937, 
    1708, 
    3488, 
    914, 
    1708, 
    2259, 
    3488, 
    3783, 
    5124, 
    3644, 
    3559, 
    2241, 
    1691, 
    3249, 
    3559, 
    2831, 
    6336, 
    2815, 
    4262, 
    3559, 
    6336, 
    4262, 
    3249, 
    3772, 
    6336, 
    2493, 
    3500, 
    2056, 
    1406, 
    2493, 
    2056, 
    5222, 
    3870, 
    6167, 
    886, 
    5222, 
    4717, 
    3601, 
    3870, 
    5222, 
    3249, 
    2831, 
    3181, 
    1691, 
    886, 
    2831, 
    2738, 
    2484, 
    736, 
    5404, 
    4334, 
    2738, 
    2159, 
    5404, 
    1572, 
    2448, 
    5303, 
    5404, 
    5303, 
    2866, 
    3217, 
    4334, 
    5303, 
    4125, 
    4334, 
    5404, 
    5303, 
    865, 
    1873, 
    5826, 
    1531, 
    1166, 
    672, 
    2237, 
    2015, 
    1685, 
    3084, 
    2237, 
    1685, 
    6022, 
    3084, 
    1685, 
    879, 
    6022, 
    1685, 
    2742, 
    3709, 
    6022, 
    5826, 
    1455, 
    865, 
    3157, 
    5873, 
    2802, 
    4151, 
    1455, 
    5826, 
    3477, 
    4363, 
    5873, 
    5051, 
    2088, 
    4151, 
    4363, 
    5051, 
    4151, 
    2708, 
    951, 
    5051, 
    879, 
    2742, 
    6022, 
    951, 
    2088, 
    5051, 
    1218, 
    822, 
    2237, 
    2119, 
    1282, 
    1978, 
    1017, 
    2912, 
    2119, 
    3906, 
    4611, 
    1266, 
    5603, 
    4366, 
    4155, 
    3240, 
    5603, 
    2900, 
    6522, 
    6189, 
    4563, 
    3240, 
    6522, 
    5603, 
    3240, 
    6189, 
    6522, 
    4744, 
    4569, 
    2698, 
    3253, 
    4916, 
    3562, 
    4611, 
    4782, 
    4857, 
    1266, 
    4611, 
    2270, 
    3906, 
    4155, 
    4782, 
    2872, 
    4620, 
    4791, 
    6295, 
    2484, 
    2900, 
    5603, 
    6295, 
    2900, 
    4155, 
    3906, 
    6295, 
    5929, 
    6053, 
    1738, 
    3824, 
    6484, 
    2479, 
    6053, 
    4510, 
    951, 
    6415, 
    6053, 
    5929, 
    2895, 
    6415, 
    5929, 
    5506, 
    6053, 
    6415, 
    5694, 
    4510, 
    6053, 
    6484, 
    5842, 
    5506, 
    2479, 
    6484, 
    5506, 
    3824, 
    4910, 
    6484, 
    4308, 
    4510, 
    5694, 
    2895, 
    5929, 
    1518, 
    5929, 
    1738, 
    2282, 
    1518, 
    5929, 
    2282, 
    2895, 
    2479, 
    6415, 
    2619, 
    2895, 
    1518, 
    2479, 
    5506, 
    6415, 
    951, 
    2708, 
    3709, 
    2742, 
    879, 
    2043, 
    2885, 
    5267, 
    2469, 
    3709, 
    2708, 
    6022, 
    2088, 
    1455, 
    4151, 
    2237, 
    822, 
    2015, 
    3084, 
    4560, 
    2237, 
    2802, 
    5873, 
    5826, 
    5694, 
    6053, 
    5506, 
    2738, 
    736, 
    1572, 
    5826, 
    1873, 
    2802, 
    1085, 
    822, 
    1218, 
    5240, 
    1866, 
    1122, 
    1004, 
    6209, 
    4465, 
    3235, 
    2473, 
    5240, 
    6212, 
    1291, 
    1192, 
    5307, 
    6212, 
    1192, 
    5307, 
    4135, 
    6212, 
    3235, 
    3874, 
    2473, 
    1982, 
    1291, 
    3874, 
    6079, 
    3344, 
    3009, 
    1866, 
    5549, 
    5282, 
    2383, 
    3344, 
    5549, 
    5307, 
    1443, 
    4135, 
    2594, 
    2838, 
    939, 
    3504, 
    3188, 
    2622, 
    5243, 
    3504, 
    3009, 
    5243, 
    3648, 
    3504, 
    3344, 
    5243, 
    3009, 
    3344, 
    1443, 
    5243, 
    2079, 
    2838, 
    3648, 
    5197, 
    2594, 
    4347, 
    939, 
    2838, 
    2079, 
    4136, 
    4347, 
    3672, 
    5549, 
    6079, 
    5282, 
    6398, 
    1166, 
    5182, 
    6191, 
    6398, 
    6079, 
    6191, 
    2158, 
    6398, 
    1932, 
    2158, 
    1085, 
    672, 
    1166, 
    2158, 
    1896, 
    5392, 
    5182, 
    735, 
    1896, 
    1166, 
    735, 
    1966, 
    2408, 
    1588, 
    754, 
    3513, 
    3584, 
    2172, 
    1588, 
    1922, 
    3584, 
    1064, 
    1922, 
    695, 
    4643, 
    1790, 
    1017, 
    754, 
    2172, 
    2328, 
    1588, 
    5405, 
    5306, 
    3485, 
    2758, 
    5405, 
    2454, 
    3123, 
    5306, 
    5405, 
    4770, 
    4468, 
    4260, 
    2654, 
    4770, 
    4228, 
    4601, 
    4468, 
    4770, 
    1790, 
    4601, 
    2654, 
    2328, 
    1343, 
    4651, 
    3166, 
    2812, 
    2454, 
    5405, 
    3166, 
    2454, 
    6546, 
    2836, 
    4260, 
    5811, 
    5947, 
    6546, 
    5947, 
    6069, 
    6491, 
    5659, 
    5811, 
    5976, 
    6413, 
    2801, 
    5491, 
    1588, 
    2328, 
    1790, 
    5290, 
    5384, 
    5726, 
    4857, 
    4689, 
    4569, 
    4916, 
    5011, 
    4744, 
    4782, 
    4689, 
    4857, 
    3906, 
    4782, 
    4611, 
    4155, 
    4366, 
    4782, 
    2043, 
    879, 
    2326, 
    2469, 
    2043, 
    899, 
    1699, 
    3542, 
    899, 
    5267, 
    2282, 
    1738, 
    3709, 
    1738, 
    951, 
    3084, 
    6022, 
    2708, 
    5267, 
    2885, 
    2282, 
    2742, 
    5267, 
    3709, 
    2742, 
    2469, 
    5267, 
    3709, 
    5267, 
    1738, 
    1282, 
    1518, 
    2282, 
    2119, 
    1518, 
    1282, 
    1790, 
    2654, 
    1017, 
    2119, 
    2912, 
    2619, 
    2469, 
    2742, 
    2043, 
    1932, 
    1085, 
    1218, 
    4363, 
    5891, 
    5051, 
    672, 
    2158, 
    1932, 
    3542, 
    2885, 
    2469, 
    5673, 
    3542, 
    1699, 
    1821, 
    5673, 
    1699, 
    1821, 
    3513, 
    5673, 
    6284, 
    1978, 
    1282, 
    5673, 
    5262, 
    3542, 
    3513, 
    754, 
    5262, 
    1341, 
    879, 
    1685, 
    2015, 
    1341, 
    1685, 
    2594, 
    5197, 
    2838, 
    822, 
    3188, 
    2015, 
    2622, 
    3009, 
    3504, 
    822, 
    2622, 
    3188, 
    3039, 
    1724, 
    2271, 
    2015, 
    3188, 
    5068, 
    939, 
    1724, 
    2594, 
    4643, 
    3584, 
    1922, 
    1821, 
    1516, 
    1064, 
    3513, 
    5262, 
    5673, 
    1017, 
    1978, 
    754, 
    3542, 
    2469, 
    899, 
    1282, 
    2885, 
    6284, 
    1282, 
    2282, 
    2885, 
    5879, 
    1789, 
    3269, 
    4870, 
    5879, 
    3269, 
    4870, 
    1699, 
    5879, 
    6266, 
    3957, 
    2797, 
    3472, 
    6507, 
    3153, 
    3689, 
    3957, 
    6266, 
    1821, 
    1699, 
    1516, 
    3584, 
    3513, 
    1064, 
    6284, 
    5262, 
    1978, 
    3542, 
    6284, 
    2885, 
    3542, 
    5262, 
    6284, 
    1064, 
    3513, 
    1821, 
    754, 
    1978, 
    5262, 
    3269, 
    1789, 
    2326, 
    2457, 
    5406, 
    3059, 
    5879, 
    1699, 
    899, 
    4698, 
    4870, 
    3269, 
    4698, 
    5406, 
    4870, 
    3575, 
    3269, 
    3672, 
    3848, 
    3575, 
    3371, 
    3039, 
    5424, 
    3371, 
    4959, 
    5099, 
    4074, 
    4806, 
    3392, 
    3059, 
    3575, 
    6112, 
    4698, 
    5668, 
    4115, 
    5099, 
    4806, 
    6112, 
    4959, 
    3848, 
    4115, 
    5668, 
    2043, 
    1789, 
    899, 
    1267, 
    5424, 
    2271, 
    4757, 
    1088, 
    797, 
    5797, 
    6447, 
    3933, 
    3575, 
    4698, 
    3269, 
    5406, 
    4806, 
    3059, 
    4870, 
    5406, 
    2457, 
    4698, 
    4806, 
    5406, 
    1699, 
    4870, 
    2457, 
    3575, 
    3848, 
    6112, 
    4959, 
    3689, 
    3392, 
    2160, 
    3957, 
    1573, 
    6266, 
    2797, 
    3153, 
    4074, 
    3957, 
    3689, 
    2160, 
    2797, 
    3957, 
    6507, 
    6266, 
    3153, 
    3392, 
    6507, 
    4603, 
    3689, 
    6266, 
    6507, 
    5616, 
    1516, 
    2457, 
    4643, 
    2172, 
    3584, 
    1088, 
    2797, 
    2160, 
    2371, 
    715, 
    1673, 
    2016, 
    1851, 
    825, 
    1102, 
    4643, 
    1851, 
    2603, 
    5458, 
    2028, 
    4597, 
    1662, 
    3385, 
    4597, 
    2222, 
    1662, 
    4397, 
    4597, 
    3385, 
    4397, 
    6136, 
    4597, 
    1190, 
    1736, 
    2222, 
    1190, 
    948, 
    1736, 
    6388, 
    1515, 
    3374, 
    2586, 
    760, 
    1596, 
    2038, 
    1384, 
    1745, 
    959, 
    2038, 
    1745, 
    3619, 
    6097, 
    3888, 
    3615, 
    3209, 
    3308, 
    4566, 
    2683, 
    1526, 
    3336, 
    4566, 
    3642, 
    4374, 
    5687, 
    4566, 
    3000, 
    4374, 
    3336, 
    4374, 
    6224, 
    5687, 
    5950, 
    3209, 
    3521, 
    6505, 
    3312, 
    2972, 
    6097, 
    3619, 
    6233, 
    2573, 
    6097, 
    2968, 
    2573, 
    3888, 
    6097, 
    2718, 
    3093, 
    3619, 
    3615, 
    2439, 
    3209, 
    6505, 
    4898, 
    3615, 
    6233, 
    6505, 
    3308, 
    6233, 
    3312, 
    6505, 
    4898, 
    2972, 
    5043, 
    2439, 
    2683, 
    3209, 
    1816, 
    1059, 
    4506, 
    5221, 
    1816, 
    4506, 
    3856, 
    5221, 
    1290, 
    2348, 
    1816, 
    5221, 
    2287, 
    3856, 
    1290, 
    4943, 
    2348, 
    1384, 
    2700, 
    4943, 
    2681, 
    5359, 
    2917, 
    3259, 
    2700, 
    5261, 
    4943, 
    2700, 
    5154, 
    5261, 
    4201, 
    4517, 
    2892, 
    4867, 
    3405, 
    3703, 
    5935, 
    4867, 
    4694, 
    2705, 
    5935, 
    4694, 
    2705, 
    3081, 
    5935, 
    3081, 
    3410, 
    5413, 
    3405, 
    2529, 
    3703, 
    3981, 
    2578, 
    3714, 
    3225, 
    3981, 
    3714, 
    872, 
    1681, 
    3981, 
    3981, 
    1681, 
    2578, 
    4107, 
    3567, 
    3841, 
    2344, 
    4107, 
    4104, 
    1374, 
    3567, 
    4107, 
    4321, 
    4107, 
    3841, 
    4106, 
    4321, 
    3841, 
    4201, 
    4104, 
    4321, 
    4292, 
    4076, 
    2718, 
    2459, 
    4404, 
    4208, 
    4190, 
    4076, 
    4292, 
    2476, 
    4190, 
    4404, 
    2476, 
    2529, 
    4190, 
    4506, 
    4627, 
    760, 
    6499, 
    1801, 
    1035, 
    2537, 
    6499, 
    6122, 
    2537, 
    2338, 
    6499, 
    5244, 
    4661, 
    2623, 
    3484, 
    4918, 
    4746, 
    3484, 
    1035, 
    4918, 
    2684, 
    4879, 
    1455, 
    2088, 
    2684, 
    1455, 
    2900, 
    2484, 
    2738, 
    4334, 
    2900, 
    2738, 
    4334, 
    5364, 
    2900, 
    3529, 
    3861, 
    3217, 
    5166, 
    3826, 
    3553, 
    3590, 
    5166, 
    3861, 
    3590, 
    5711, 
    5166, 
    4738, 
    4910, 
    4091, 
    3824, 
    3342, 
    3647, 
    5016, 
    3342, 
    3006, 
    4002, 
    5016, 
    2498, 
    4863, 
    3342, 
    5016, 
    3449, 
    4863, 
    3737, 
    4692, 
    3647, 
    4863, 
    4091, 
    3824, 
    3647, 
    5708, 
    4305, 
    6025, 
    3403, 
    5708, 
    3701, 
    3403, 
    5128, 
    5708, 
    4305, 
    4563, 
    4738, 
    3824, 
    2479, 
    3342, 
    6025, 
    4091, 
    3647, 
    3701, 
    6025, 
    3647, 
    3701, 
    5708, 
    6025, 
    4510, 
    2684, 
    2088, 
    1738, 
    6053, 
    951, 
    4308, 
    2684, 
    4510, 
    6484, 
    4910, 
    6367, 
    4092, 
    4879, 
    4308, 
    6367, 
    4910, 
    4738, 
    4308, 
    5842, 
    4092, 
    5694, 
    5506, 
    5842, 
    5711, 
    3590, 
    3283, 
    5966, 
    5711, 
    3283, 
    5029, 
    5166, 
    5711, 
    4092, 
    5029, 
    4879, 
    3826, 
    5166, 
    5029, 
    6189, 
    4738, 
    4563, 
    4092, 
    6367, 
    3826, 
    6367, 
    4738, 
    6082, 
    4308, 
    5694, 
    5842, 
    3824, 
    4091, 
    4910, 
    3553, 
    5266, 
    5166, 
    5698, 
    4366, 
    4563, 
    4689, 
    5698, 
    4508, 
    4689, 
    4366, 
    5698, 
    5128, 
    4689, 
    4508, 
    5708, 
    5128, 
    4508, 
    3074, 
    4569, 
    5128, 
    4569, 
    4744, 
    4857, 
    2484, 
    6295, 
    3906, 
    6082, 
    3553, 
    3826, 
    4508, 
    4563, 
    4305, 
    4366, 
    5603, 
    6522, 
    2159, 
    2448, 
    5404, 
    2159, 
    1086, 
    2448, 
    3165, 
    2159, 
    1572, 
    736, 
    5325, 
    1572, 
    4918, 
    2130, 
    4661, 
    6122, 
    3484, 
    3165, 
    5325, 
    6122, 
    3165, 
    5325, 
    2537, 
    6122, 
    1035, 
    2130, 
    4918, 
    4398, 
    1838, 
    3456, 
    4746, 
    4985, 
    2159, 
    3613, 
    2815, 
    3169, 
    4212, 
    3883, 
    3613, 
    4661, 
    4212, 
    2623, 
    680, 
    3883, 
    4212, 
    680, 
    1937, 
    3883, 
    4426, 
    5209, 
    680, 
    3772, 
    2493, 
    1406, 
    3169, 
    3772, 
    1406, 
    3169, 
    2815, 
    3772, 
    1838, 
    3010, 
    3169, 
    4262, 
    2241, 
    3559, 
    5124, 
    2615, 
    3644, 
    4269, 
    5124, 
    4043, 
    4162, 
    2615, 
    5124, 
    4269, 
    4478, 
    5124, 
    3339, 
    2796, 
    4162, 
    1617, 
    3152, 
    786, 
    6077, 
    4948, 
    2796, 
    1134, 
    2848, 
    2187, 
    4398, 
    2448, 
    1086, 
    3772, 
    2815, 
    6336, 
    1838, 
    3169, 
    2360, 
    3010, 
    2623, 
    3613, 
    5380, 
    2615, 
    4948, 
    1406, 
    5380, 
    4721, 
    1406, 
    2056, 
    5380, 
    3339, 
    786, 
    3152, 
    4721, 
    2360, 
    1406, 
    4948, 
    4721, 
    5380, 
    3132, 
    3456, 
    4721, 
    3918, 
    4165, 
    2769, 
    3456, 
    2360, 
    4721, 
    4165, 
    4186, 
    5776, 
    1838, 
    2360, 
    3456, 
    4162, 
    2796, 
    2615, 
    786, 
    3339, 
    1996, 
    3152, 
    2796, 
    3339, 
    2187, 
    5276, 
    1617, 
    5276, 
    3197, 
    5176, 
    5766, 
    2487, 
    2902, 
    5126, 
    4836, 
    2660, 
    3377, 
    5241, 
    3044, 
    3611, 
    4836, 
    5126, 
    2964, 
    3305, 
    2569, 
    1617, 
    786, 
    4836, 
    786, 
    1996, 
    2660, 
    4948, 
    3132, 
    4721, 
    2796, 
    4948, 
    2615, 
    2769, 
    3132, 
    4948, 
    6188, 
    1296, 
    4813, 
    3923, 
    2210, 
    1169, 
    5198, 
    4049, 
    3923, 
    2627, 
    5198, 
    3923, 
    1751, 
    1044, 
    2135, 
    2057, 
    1751, 
    1408, 
    3004, 
    3903, 
    1408, 
    907, 
    1751, 
    2057, 
    907, 
    967, 
    1751, 
    4664, 
    1169, 
    1898, 
    1703, 
    4664, 
    1898, 
    2627, 
    3923, 
    4664, 
    4839, 
    2627, 
    4664, 
    907, 
    4839, 
    1703, 
    3014, 
    2627, 
    4839, 
    2057, 
    3014, 
    907, 
    5198, 
    2617, 
    3788, 
    2057, 
    3903, 
    3014, 
    2057, 
    1408, 
    3903, 
    3014, 
    5198, 
    2627, 
    4664, 
    3923, 
    1169, 
    1649, 
    1420, 
    2210, 
    5198, 
    3903, 
    2617, 
    4049, 
    5198, 
    3788, 
    3014, 
    3903, 
    5198, 
    1851, 
    2371, 
    825, 
    4940, 
    1811, 
    917, 
    1420, 
    4940, 
    2210, 
    1420, 
    863, 
    4940, 
    2371, 
    1673, 
    1420, 
    1649, 
    2371, 
    1420, 
    1851, 
    715, 
    2371, 
    863, 
    1811, 
    4940, 
    917, 
    167, 
    1898, 
    1703, 
    165, 
    967, 
    2292, 
    807, 
    1300, 
    972, 
    1764, 
    1757, 
    5484, 
    2817, 
    3170, 
    1757, 
    1764, 
    1634, 
    4264, 
    2599, 
    5052, 
    4471, 
    4264, 
    2794, 
    4562, 
    4471, 
    3151, 
    4168, 
    4562, 
    3151, 
    1585, 
    2170, 
    4830, 
    5534, 
    2853, 
    6119, 
    4471, 
    5534, 
    6119, 
    5572, 
    5777, 
    2599, 
    6119, 
    5572, 
    2599, 
    5249, 
    5299, 
    6432, 
    5963, 
    5200, 
    5553, 
    6245, 
    5963, 
    5553, 
    5677, 
    5299, 
    5963, 
    5777, 
    6432, 
    5677, 
    5998, 
    5586, 
    5861, 
    5249, 
    5519, 
    5299, 
    6163, 
    2433, 
    2853, 
    6098, 
    5486, 
    5755, 
    5998, 
    5861, 
    5849, 
    3345, 
    5998, 
    3649, 
    3345, 
    5586, 
    5998, 
    5861, 
    6458, 
    5849, 
    6396, 
    6023, 
    6142, 
    6244, 
    6404, 
    6142, 
    6264, 
    6163, 
    6396, 
    6501, 
    6163, 
    6264, 
    6501, 
    2433, 
    6163, 
    6445, 
    6408, 
    5632, 
    5486, 
    6551, 
    5755, 
    6331, 
    6403, 
    6409, 
    6331, 
    5679, 
    6264, 
    6386, 
    4663, 
    5946, 
    6023, 
    6386, 
    6142, 
    6023, 
    3202, 
    6386, 
    6501, 
    5249, 
    2433, 
    5679, 
    6501, 
    6264, 
    5519, 
    5249, 
    6501, 
    2853, 
    3202, 
    6023, 
    5519, 
    5720, 
    5299, 
    2633, 
    6261, 
    5553, 
    927, 
    4168, 
    1279, 
    2817, 
    6035, 
    5052, 
    1165, 
    1891, 
    5916, 
    4284, 
    4492, 
    2667, 
    5792, 
    5632, 
    5752, 
    5894, 
    5792, 
    4379, 
    6561, 
    6445, 
    5632, 
    5894, 
    6561, 
    5792, 
    5894, 
    5755, 
    6561, 
    3919, 
    5985, 
    6098, 
    6428, 
    6318, 
    5552, 
    5730, 
    6429, 
    5552, 
    6553, 
    6547, 
    6537, 
    6428, 
    6553, 
    6506, 
    6410, 
    6547, 
    6553, 
    6509, 
    6410, 
    5670, 
    5474, 
    6509, 
    5670, 
    6408, 
    6547, 
    6509, 
    6408, 
    6508, 
    6547, 
    5474, 
    6408, 
    6509, 
    6403, 
    6396, 
    6404, 
    6403, 
    6264, 
    6396, 
    6404, 
    6537, 
    6403, 
    6551, 
    5486, 
    5679, 
    6409, 
    6551, 
    6331, 
    6409, 
    6508, 
    6563, 
    6429, 
    5954, 
    5818, 
    5552, 
    6429, 
    6428, 
    5730, 
    5954, 
    6429, 
    5892, 
    6043, 
    4065, 
    5894, 
    4379, 
    4166, 
    6098, 
    5894, 
    4166, 
    3919, 
    6098, 
    4166, 
    5985, 
    5486, 
    6098, 
    5755, 
    6563, 
    6561, 
    6547, 
    6410, 
    6509, 
    6537, 
    6547, 
    6508, 
    6537, 
    6404, 
    6553, 
    5792, 
    4572, 
    4379, 
    5587, 
    5752, 
    5632, 
    6552, 
    6435, 
    6012, 
    5752, 
    6552, 
    6469, 
    5587, 
    6435, 
    6552, 
    6271, 
    6056, 
    3934, 
    3362, 
    6271, 
    3663, 
    5607, 
    6056, 
    6271, 
    5059, 
    6128, 
    5192, 
    6128, 
    5741, 
    6056, 
    5783, 
    5917, 
    5741, 
    3804, 
    3525, 
    5567, 
    4275, 
    3546, 
    4572, 
    4663, 
    3516, 
    3796, 
    915, 
    2883, 
    2064, 
    3362, 
    2367, 
    1413, 
    683, 
    1256, 
    1585, 
    3212, 
    4852, 
    2862, 
    5442, 
    1565, 
    5310, 
    2152, 
    780, 
    889, 
    5310, 
    1565, 
    2152, 
    2369, 
    5310, 
    1417, 
    2369, 
    5442, 
    5310, 
    2064, 
    2443, 
    1417, 
    5442, 
    725, 
    1565, 
    1848, 
    5442, 
    2369, 
    1848, 
    4512, 
    5442, 
    725, 
    1614, 
    1565, 
    1993, 
    807, 
    821, 
    6245, 
    3170, 
    5677, 
    783, 
    4741, 
    1993, 
    1723, 
    2270, 
    5011, 
    6380, 
    5947, 
    6358, 
    5706, 
    5975, 
    5501, 
    3485, 
    6069, 
    5975, 
    5306, 
    3449, 
    5884, 
    3166, 
    5405, 
    3485, 
    3123, 
    3449, 
    5306, 
    4002, 
    3737, 
    5016, 
    3485, 
    5306, 
    3186, 
    5508, 
    3403, 
    3701, 
    4692, 
    5508, 
    3701, 
    3123, 
    2758, 
    5508, 
    3074, 
    3403, 
    2758, 
    5884, 
    3737, 
    5502, 
    2619, 
    2498, 
    3006, 
    2895, 
    2619, 
    3006, 
    1518, 
    2119, 
    2619, 
    1790, 
    2328, 
    4601, 
    1872, 
    1003, 
    1014, 
    4676, 
    6181, 
    1014, 
    1515, 
    4815, 
    1872, 
    1779, 
    1003, 
    5336, 
    4030, 
    2417, 
    1452, 
    4073, 
    1910, 
    1190, 
    4714, 
    2382, 
    3754, 
    1910, 
    4030, 
    1190, 
    2111, 
    1872, 
    4815, 
    1501, 
    6007, 
    2111, 
    1003, 
    1872, 
    2111, 
    6388, 
    6049, 
    1921, 
    1515, 
    6388, 
    1452, 
    3374, 
    6049, 
    6388, 
    6181, 
    4676, 
    5633, 
    1872, 
    6181, 
    1515, 
    1872, 
    1014, 
    6181, 
    3041, 
    5881, 
    6049, 
    4687, 
    3011, 
    3345, 
    4507, 
    6525, 
    4687, 
    4676, 
    3011, 
    4687, 
    3374, 
    6181, 
    5633, 
    1014, 
    2624, 
    4676, 
    5631, 
    2901, 
    3241, 
    5881, 
    5631, 
    3241, 
    2657, 
    4390, 
    5631, 
    4815, 
    1515, 
    1452, 
    2417, 
    4815, 
    1452, 
    1501, 
    2111, 
    4815, 
    5792, 
    5752, 
    4572, 
    5783, 
    6435, 
    5474, 
    6469, 
    4275, 
    4572, 
    5587, 
    6552, 
    5752, 
    4919, 
    4275, 
    6469, 
    6012, 
    5059, 
    4919, 
    6469, 
    6552, 
    4919, 
    6128, 
    5607, 
    5192, 
    5584, 
    6128, 
    6012, 
    5584, 
    5741, 
    6128, 
    5670, 
    5783, 
    5474, 
    6271, 
    3934, 
    3663, 
    6128, 
    6056, 
    5607, 
    6534, 
    3934, 
    6056, 
    5741, 
    6534, 
    6056, 
    5741, 
    5567, 
    6534, 
    5783, 
    5741, 
    5584, 
    6435, 
    5783, 
    5584, 
    5670, 
    5818, 
    5917, 
    5567, 
    3525, 
    6534, 
    2655, 
    4275, 
    2890, 
    3804, 
    5567, 
    5892, 
    3546, 
    4379, 
    4572, 
    2853, 
    6023, 
    6163, 
    5587, 
    5632, 
    5474, 
    5755, 
    5894, 
    6098, 
    3822, 
    4166, 
    4379, 
    5985, 
    3649, 
    5998, 
    5486, 
    5985, 
    5849, 
    3919, 
    3649, 
    5985, 
    4865, 
    5992, 
    3960, 
    4284, 
    4083, 
    4065, 
    2667, 
    4773, 
    4083, 
    3384, 
    848, 
    1662, 
    4555, 
    3384, 
    1662, 
    1278, 
    4621, 
    3384, 
    2281, 
    1672, 
    1278, 
    4555, 
    1736, 
    2281, 
    5636, 
    5793, 
    3554, 
    862, 
    2036, 
    1977, 
    750, 
    4574, 
    1977, 
    4574, 
    1364, 
    2028, 
    1584, 
    4574, 
    750, 
    1584, 
    5354, 
    4574, 
    1374, 
    1584, 
    750, 
    5500, 
    4650, 
    1801, 
    5354, 
    5500, 
    1801, 
    5354, 
    2169, 
    5500, 
    2338, 
    2537, 
    1364, 
    2088, 
    951, 
    4510, 
    1472, 
    5091, 
    139, 
    4276, 
    1261, 
    3155, 
    4469, 
    1757, 
    2292, 
    4261, 
    4469, 
    4247, 
    5111, 
    972, 
    1757, 
    4261, 
    5111, 
    4469, 
    4261, 
    5329, 
    5111, 
    4017, 
    4261, 
    4247, 
    5329, 
    4276, 
    4485, 
    4036, 
    5329, 
    4261, 
    4036, 
    5417, 
    5329, 
    2560, 
    1079, 
    2156, 
    1568, 
    2560, 
    2156, 
    4829, 
    932, 
    6129, 
    6038, 
    4829, 
    2941, 
    1834, 
    6038, 
    2941, 
    1079, 
    2560, 
    6038, 
    1720, 
    932, 
    4829, 
    4469, 
    5111, 
    1757, 
    2783, 
    4036, 
    4017, 
    5417, 
    1447, 
    4276, 
    3771, 
    5417, 
    4036, 
    3771, 
    1720, 
    5417, 
    1720, 
    4829, 
    2560, 
    1938, 
    2156, 
    1224, 
    6050, 
    2626, 
    3013, 
    4485, 
    3155, 
    1891, 
    5417, 
    4276, 
    5329, 
    1447, 
    1261, 
    4276, 
    4455, 
    2292, 
    1300, 
    3771, 
    4036, 
    2783, 
    4469, 
    2292, 
    4455, 
    1987, 
    1300, 
    807, 
    1993, 
    4741, 
    807, 
    4255, 
    1605, 
    2179, 
    3027, 
    3787, 
    2641, 
    3476, 
    6140, 
    3764, 
    4016, 
    3751, 
    3908, 
    6003, 
    4016, 
    2561, 
    1861, 
    6003, 
    2561, 
    1271, 
    3348, 
    6003, 
    6527, 
    5639, 
    3751, 
    6003, 
    6527, 
    4016, 
    6003, 
    3348, 
    6527, 
    1435, 
    1728, 
    5627, 
    5782, 
    3464, 
    5639, 
    3013, 
    5782, 
    5639, 
    2626, 
    3111, 
    5782, 
    932, 
    1720, 
    3771, 
    5365, 
    770, 
    1605, 
    5447, 
    5224, 
    5365, 
    5093, 
    5245, 
    5224, 
    5959, 
    4819, 
    2536, 
    4979, 
    5649, 
    4826, 
    6473, 
    1337, 
    151, 
    6221, 
    5649, 
    5334, 
    4979, 
    894, 
    5802, 
    5802, 
    4972, 
    5334, 
    4979, 
    5802, 
    5649, 
    6473, 
    1401, 
    4972, 
    1337, 
    6473, 
    5802, 
    151, 
    1401, 
    6473, 
    1401, 
    2357, 
    4972, 
    3329, 
    696, 
    1946, 
    4365, 
    2991, 
    2601, 
    325, 
    4365, 
    2601, 
    324, 
    902, 
    4365, 
    902, 
    696, 
    2991, 
    1228, 
    3295, 
    4926, 
    1700, 
    2251, 
    6288, 
    4421, 
    2104, 
    3247, 
    1236, 
    4421, 
    3247, 
    1946, 
    696, 
    4421, 
    5063, 
    4926, 
    3602, 
    3871, 
    5063, 
    3602, 
    902, 
    4577, 
    5063, 
    5922, 
    5737, 
    3696, 
    3963, 
    5922, 
    3696, 
    4313, 
    4096, 
    6489, 
    1539, 
    5260, 
    4096, 
    2133, 
    4762, 
    5260, 
    5922, 
    6489, 
    5737, 
    5488, 
    2691, 
    3963, 
    2468, 
    5488, 
    3963, 
    2884, 
    1766, 
    5488, 
    3871, 
    1484, 
    5063, 
    5759, 
    3153, 
    2797, 
    4930, 
    5759, 
    4757, 
    6535, 
    5069, 
    5931, 
    6470, 
    5797, 
    4174, 
    4930, 
    5069, 
    6535, 
    5069, 
    5837, 
    5931, 
    3431, 
    5069, 
    4930, 
    2731, 
    5296, 
    5837, 
    3933, 
    3760, 
    4174, 
    3760, 
    3472, 
    4174, 
    4025, 
    3760, 
    3933, 
    5955, 
    4251, 
    4025, 
    3361, 
    5955, 
    3662, 
    3361, 
    715, 
    5955, 
    4771, 
    3059, 
    4603, 
    3760, 
    4771, 
    4603, 
    4483, 
    5616, 
    4771, 
    4251, 
    4483, 
    4025, 
    1922, 
    1064, 
    6440, 
    4025, 
    4483, 
    4771, 
    4603, 
    3059, 
    3392, 
    5627, 
    1728, 
    3142, 
    6050, 
    5627, 
    3142, 
    3348, 
    1435, 
    5627, 
    783, 
    1616, 
    2317, 
    3111, 
    2744, 
    6140, 
    3464, 
    5782, 
    3141, 
    5428, 
    2783, 
    4017, 
    4785, 
    2179, 
    1605, 
    5268, 
    4785, 
    1605, 
    1779, 
    5336, 
    4785, 
    5190, 
    1865, 
    2382, 
    5190, 
    4481, 
    1865, 
    3533, 
    5290, 
    3811, 
    6067, 
    5726, 
    2641, 
    4481, 
    6067, 
    4273, 
    5290, 
    5726, 
    6067, 
    3811, 
    5290, 
    5190, 
    3533, 
    3222, 
    5384, 
    5187, 
    2179, 
    1120, 
    4273, 
    5187, 
    4481, 
    4273, 
    5055, 
    5187, 
    6597, 
    163, 
    5134, 
    165, 
    6597, 
    967, 
    165, 
    164, 
    6597, 
    4499, 
    2115, 
    3656, 
    4582, 
    5129, 
    1601, 
    4755, 
    6243, 
    4582, 
    5928, 
    4826, 
    4647, 
    4837, 
    5928, 
    4983, 
    4837, 
    4979, 
    5928, 
    3656, 
    1510, 
    2031, 
    155, 
    2205, 
    4499, 
    1010, 
    1231, 
    2115, 
    5091, 
    3155, 
    1261, 
    139, 
    5091, 
    729, 
    1472, 
    3155, 
    5091, 
    4168, 
    3926, 
    1279, 
    5916, 
    2786, 
    3926, 
    2670, 
    6146, 
    2786, 
    1891, 
    1472, 
    2670, 
    138, 
    1431, 
    139, 
    137, 
    1279, 
    1431, 
    4168, 
    751, 
    4562, 
    3926, 
    4168, 
    3151, 
    927, 
    751, 
    4168, 
    5245, 
    1300, 
    1987, 
    5224, 
    5245, 
    1987, 
    5093, 
    5345, 
    5245, 
    5345, 
    4455, 
    5245, 
    4247, 
    4469, 
    4455, 
    3111, 
    2626, 
    5428, 
    4017, 
    4036, 
    4261, 
    5417, 
    1720, 
    1447, 
    3142, 
    3771, 
    2783, 
    3142, 
    932, 
    3771, 
    1757, 
    1634, 
    2292, 
    1165, 
    1764, 
    972, 
    1634, 
    807, 
    2292, 
    2016, 
    1343, 
    1102, 
    4228, 
    4770, 
    4939, 
    6263, 
    6407, 
    6352, 
    4173, 
    3932, 
    6294, 
    6491, 
    6546, 
    5947, 
    4468, 
    6124, 
    4260, 
    5655, 
    5659, 
    5976, 
    6162, 
    5942, 
    6045, 
    3004, 
    5808, 
    2617, 
    6066, 
    4756, 
    4583, 
    5919, 
    6066, 
    4583, 
    5942, 
    5482, 
    6066, 
    4737, 
    2210, 
    3923, 
    4482, 
    4737, 
    4274, 
    1649, 
    2210, 
    4737, 
    4274, 
    3923, 
    4049, 
    4274, 
    4737, 
    3923, 
    3332, 
    1577, 
    743, 
    3638, 
    3332, 
    2561, 
    6412, 
    3660, 
    3932, 
    5491, 
    6412, 
    3932, 
    5491, 
    3190, 
    6412, 
    5520, 
    3660, 
    3359, 
    3027, 
    5606, 
    5648, 
    6294, 
    5623, 
    5785, 
    4173, 
    6294, 
    5785, 
    5836, 
    5691, 
    6294, 
    3660, 
    5836, 
    3932, 
    5691, 
    5623, 
    6294, 
    6308, 
    5691, 
    5520, 
    5648, 
    6308, 
    5520, 
    5801, 
    5706, 
    6308, 
    5501, 
    6340, 
    5691, 
    5520, 
    5836, 
    3660, 
    6478, 
    6357, 
    6453, 
    6162, 
    6478, 
    6263, 
    6356, 
    6548, 
    6478, 
    6357, 
    5811, 
    5659, 
    6453, 
    6357, 
    5659, 
    6477, 
    6340, 
    6380, 
    6358, 
    6548, 
    6380, 
    6356, 
    6443, 
    6477, 
    6045, 
    6356, 
    6162, 
    6358, 
    5947, 
    5811, 
    6548, 
    6477, 
    6380, 
    6478, 
    6548, 
    6357, 
    6356, 
    6477, 
    6548, 
    6380, 
    5975, 
    6069, 
    6357, 
    6548, 
    6358, 
    6340, 
    5501, 
    6380, 
    6069, 
    5947, 
    6380, 
    3186, 
    6069, 
    3485, 
    3186, 
    2836, 
    6491, 
    6069, 
    3186, 
    6491, 
    6546, 
    6491, 
    2836, 
    5976, 
    6546, 
    4260, 
    5976, 
    5811, 
    6546, 
    5691, 
    5836, 
    5520, 
    2840, 
    4929, 
    5482, 
    4385, 
    5555, 
    4173, 
    5491, 
    2801, 
    3190, 
    4173, 
    6542, 
    3932, 
    6542, 
    5555, 
    6413, 
    5491, 
    6542, 
    6413, 
    4173, 
    5555, 
    6542, 
    2561, 
    4016, 
    3638, 
    6412, 
    3190, 
    3660, 
    6413, 
    3908, 
    2801, 
    3932, 
    6542, 
    5491, 
    5555, 
    3908, 
    6413, 
    4583, 
    6337, 
    4385, 
    3638, 
    3908, 
    5555, 
    4568, 
    4049, 
    3788, 
    6352, 
    5808, 
    5942, 
    6330, 
    6407, 
    6263, 
    2617, 
    5808, 
    6352, 
    5690, 
    6124, 
    4651, 
    6204, 
    5659, 
    5655, 
    4568, 
    6204, 
    4743, 
    6478, 
    6162, 
    6356, 
    6453, 
    6263, 
    6478, 
    6204, 
    6453, 
    5659, 
    6330, 
    6263, 
    6453, 
    4568, 
    6330, 
    6204, 
    4568, 
    3788, 
    6330, 
    6407, 
    3788, 
    2617, 
    6352, 
    6407, 
    2617, 
    6330, 
    3788, 
    6407, 
    5976, 
    4260, 
    6124, 
    5502, 
    4939, 
    2836, 
    4915, 
    825, 
    4482, 
    6520, 
    4756, 
    5551, 
    6337, 
    6520, 
    5551, 
    4583, 
    4756, 
    6520, 
    2721, 
    4582, 
    765, 
    6243, 
    4755, 
    6051, 
    4837, 
    6243, 
    6051, 
    4983, 
    5129, 
    6243, 
    5428, 
    5345, 
    2744, 
    2783, 
    5428, 
    2626, 
    4017, 
    4247, 
    5428, 
    5365, 
    4255, 
    4029, 
    770, 
    5365, 
    5224, 
    1605, 
    4255, 
    5365, 
    3348, 
    3013, 
    6527, 
    1435, 
    3348, 
    1271, 
    5639, 
    3464, 
    3751, 
    3787, 
    3027, 
    3359, 
    3764, 
    3787, 
    3506, 
    3764, 
    4029, 
    4912, 
    5190, 
    5290, 
    6067, 
    5055, 
    2641, 
    4912, 
    2179, 
    5187, 
    4255, 
    1120, 
    1865, 
    4481, 
    5801, 
    6308, 
    5648, 
    3004, 
    5482, 
    5808, 
    3190, 
    3506, 
    3660, 
    3156, 
    3190, 
    2801, 
    5975, 
    5706, 
    3166, 
    3156, 
    3476, 
    3190, 
    5801, 
    5769, 
    5460, 
    3359, 
    3027, 
    5648, 
    3027, 
    2641, 
    5606, 
    5706, 
    2812, 
    3166, 
    3485, 
    5975, 
    3166, 
    5501, 
    5691, 
    6308, 
    3506, 
    3476, 
    3764, 
    3660, 
    3506, 
    3359, 
    3190, 
    3476, 
    3506, 
    3464, 
    3156, 
    2801, 
    3141, 
    3476, 
    3156, 
    3464, 
    3141, 
    3156, 
    3751, 
    3464, 
    2801, 
    3908, 
    3751, 
    2801, 
    5782, 
    3013, 
    2626, 
    4016, 
    6527, 
    3751, 
    6527, 
    3013, 
    5639, 
    5782, 
    3111, 
    3141, 
    3506, 
    3787, 
    3359, 
    6140, 
    3476, 
    3141, 
    3111, 
    6140, 
    3141, 
    2744, 
    5447, 
    6140, 
    3764, 
    6140, 
    5447, 
    5726, 
    5384, 
    5769, 
    2641, 
    5726, 
    5606, 
    2641, 
    4273, 
    6067, 
    5405, 
    2758, 
    3123, 
    4385, 
    6337, 
    5555, 
    5836, 
    6294, 
    3932, 
    5785, 
    4385, 
    4173, 
    6340, 
    6477, 
    5623, 
    5919, 
    4385, 
    5785, 
    5919, 
    4583, 
    4385, 
    6443, 
    6356, 
    6045, 
    5623, 
    6443, 
    5785, 
    5623, 
    6477, 
    6443, 
    6066, 
    5482, 
    4756, 
    6045, 
    5942, 
    6066, 
    5785, 
    6443, 
    5919, 
    6162, 
    6352, 
    5942, 
    5919, 
    6443, 
    6045, 
    6453, 
    6204, 
    6330, 
    5808, 
    5482, 
    5942, 
    5919, 
    6045, 
    6066, 
    2840, 
    5482, 
    3004, 
    4929, 
    4756, 
    5482, 
    1841, 
    4929, 
    2840, 
    1841, 
    765, 
    5681, 
    5551, 
    5681, 
    1601, 
    5681, 
    4929, 
    1841, 
    1601, 
    5681, 
    765, 
    5551, 
    4756, 
    5681, 
    5681, 
    4756, 
    4929, 
    3332, 
    5551, 
    1577, 
    3332, 
    3638, 
    6337, 
    2617, 
    3903, 
    3004, 
    743, 
    1861, 
    2561, 
    2422, 
    690, 
    4967, 
    2031, 
    1510, 
    2422, 
    1211, 
    2031, 
    857, 
    3656, 
    2115, 
    1510, 
    905, 
    3656, 
    2031, 
    905, 
    155, 
    3656, 
    1941, 
    690, 
    2422, 
    1231, 
    1941, 
    1510, 
    4582, 
    1601, 
    765, 
    4755, 
    4582, 
    2721, 
    1941, 
    4755, 
    2721, 
    6051, 
    1010, 
    1694, 
    4983, 
    6243, 
    4837, 
    1231, 
    1010, 
    6051, 
    4979, 
    1694, 
    894, 
    4647, 
    5179, 
    5928, 
    4755, 
    1231, 
    6051, 
    1694, 
    4837, 
    6051, 
    3810, 
    3768, 
    1694, 
    5179, 
    1861, 
    743, 
    5179, 
    4647, 
    1861, 
    5129, 
    5179, 
    743, 
    5129, 
    4983, 
    5179, 
    4979, 
    4826, 
    5928, 
    1694, 
    4979, 
    4837, 
    894, 
    1337, 
    5802, 
    5334, 
    5649, 
    5802, 
    4819, 
    5334, 
    4972, 
    2721, 
    690, 
    1941, 
    1231, 
    4755, 
    1941, 
    6188, 
    1841, 
    1296, 
    690, 
    6188, 
    4813, 
    765, 
    1841, 
    6188, 
    2381, 
    627, 
    315, 
    4762, 
    5561, 
    5260, 
    316, 
    627, 
    1183, 
    784, 
    315, 
    314, 
    2401, 
    3509, 
    314, 
    4257, 
    3462, 
    3749, 
    1154, 
    4257, 
    3790, 
    2199, 
    1636, 
    4257, 
    1157, 
    2199, 
    1154, 
    3749, 
    2293, 
    1758, 
    3509, 
    5729, 
    3863, 
    5025, 
    4700, 
    4873, 
    3462, 
    5025, 
    4873, 
    3462, 
    809, 
    5025, 
    1636, 
    3462, 
    4257, 
    1636, 
    809, 
    3462, 
    4873, 
    4528, 
    1988, 
    3749, 
    4873, 
    1302, 
    3749, 
    3462, 
    4873, 
    814, 
    2007, 
    809, 
    4528, 
    6017, 
    2544, 
    2301, 
    936, 
    2077, 
    4297, 
    1765, 
    1302, 
    1988, 
    4297, 
    1302, 
    983, 
    1765, 
    4297, 
    983, 
    1722, 
    1765, 
    2077, 
    840, 
    1655, 
    1311, 
    2077, 
    1440, 
    1311, 
    2301, 
    2077, 
    2077, 
    936, 
    840, 
    1758, 
    1311, 
    973, 
    1758, 
    2293, 
    2301, 
    1483, 
    1966, 
    1265, 
    5241, 
    5126, 
    3044, 
    5145, 
    5241, 
    3377, 
    3881, 
    5126, 
    5241, 
    3881, 
    3611, 
    5126, 
    5241, 
    4138, 
    3881, 
    3676, 
    5145, 
    3377, 
    3676, 
    2334, 
    5145, 
    5233, 
    1028, 
    2125, 
    5419, 
    5233, 
    4759, 
    4587, 
    5419, 
    4759, 
    2569, 
    3611, 
    5419, 
    4138, 
    1028, 
    5233, 
    5241, 
    5145, 
    4138, 
    1795, 
    1028, 
    4138, 
    2569, 
    3305, 
    3611, 
    3305, 
    4836, 
    3611, 
    1996, 
    1313, 
    2829, 
    1358, 
    2269, 
    2334, 
    6047, 
    2902, 
    3243, 
    4759, 
    5233, 
    2125, 
    2660, 
    2829, 
    3044, 
    2829, 
    2487, 
    3044, 
    1996, 
    2829, 
    2660, 
    1313, 
    698, 
    4472, 
    1358, 
    3676, 
    3781, 
    4266, 
    2902, 
    2487, 
    5311, 
    3696, 
    3401, 
    2902, 
    4311, 
    3243, 
    2468, 
    3696, 
    4311, 
    936, 
    2022, 
    840, 
    936, 
    1722, 
    2022, 
    3611, 
    3881, 
    5419, 
    2269, 
    1265, 
    2334, 
    1265, 
    1028, 
    1795, 
    983, 
    4682, 
    2103, 
    4615, 
    3289, 
    1607, 
    5535, 
    4615, 
    2180, 
    2606, 
    5535, 
    2180, 
    2606, 
    5392, 
    5535, 
    2408, 
    1483, 
    4615, 
    2103, 
    1483, 
    1265, 
    2269, 
    2103, 
    1265, 
    1795, 
    2334, 
    1265, 
    1722, 
    983, 
    2269, 
    4682, 
    1988, 
    772, 
    2103, 
    4682, 
    3289, 
    983, 
    4297, 
    4682, 
    5392, 
    4615, 
    5535, 
    4615, 
    1607, 
    2180, 
    2103, 
    3289, 
    1483, 
    772, 
    1607, 
    3289, 
    2949, 
    1332, 
    2318, 
    1781, 
    3086, 
    2318, 
    6017, 
    4528, 
    4700, 
    3413, 
    2180, 
    1607, 
    2318, 
    3086, 
    2949, 
    1781, 
    1004, 
    4465, 
    772, 
    1988, 
    4528, 
    735, 
    1166, 
    1531, 
    1311, 
    1440, 
    973, 
    1722, 
    2269, 
    1358, 
    4472, 
    2829, 
    1313, 
    1766, 
    4472, 
    698, 
    4266, 
    2829, 
    4472, 
    2334, 
    1795, 
    5145, 
    4478, 
    3339, 
    4162, 
    4472, 
    2884, 
    4266, 
    3644, 
    5380, 
    2056, 
    3644, 
    2615, 
    5380, 
    900, 
    3644, 
    2056, 
    4269, 
    2820, 
    698, 
    4478, 
    4162, 
    5124, 
    1313, 
    4478, 
    4269, 
    1996, 
    3339, 
    4478, 
    6288, 
    3173, 
    2820, 
    3783, 
    6288, 
    4043, 
    3783, 
    1700, 
    6288, 
    900, 
    3783, 
    3644, 
    900, 
    1700, 
    3783, 
    5276, 
    5176, 
    3152, 
    2848, 
    5276, 
    2187, 
    2848, 
    3197, 
    5276, 
    2381, 
    315, 
    784, 
    313, 
    2401, 
    314, 
    310, 
    1157, 
    1154, 
    6359, 
    865, 
    2942, 
    2964, 
    4388, 
    1134, 
    4560, 
    1932, 
    1218, 
    5891, 
    4363, 
    4560, 
    3084, 
    5891, 
    4560, 
    3084, 
    2708, 
    5891, 
    3974, 
    1531, 
    672, 
    3157, 
    3974, 
    3477, 
    5397, 
    2802, 
    4388, 
    5873, 
    4151, 
    5826, 
    3477, 
    5873, 
    3157, 
    4363, 
    4151, 
    5873, 
    4560, 
    4363, 
    3477, 
    1932, 
    4560, 
    3477, 
    1218, 
    2237, 
    4560, 
    5891, 
    2708, 
    5051, 
    5397, 
    4388, 
    4587, 
    1134, 
    4388, 
    1873, 
    672, 
    1932, 
    3477, 
    1457, 
    5027, 
    5911, 
    4570, 
    177, 
    4745, 
    3099, 
    6310, 
    1529, 
    6310, 
    4896, 
    2767, 
    1529, 
    6310, 
    1132, 
    3099, 
    6315, 
    6310, 
    6315, 
    4896, 
    6310, 
    3427, 
    6315, 
    3099, 
    3427, 
    3984, 
    6315, 
    6073, 
    3130, 
    4896, 
    5246, 
    6073, 
    4896, 
    5246, 
    5516, 
    6073, 
    6226, 
    3742, 
    5516, 
    752, 
    6226, 
    5516, 
    919, 
    1280, 
    6226, 
    4298, 
    6524, 
    3398, 
    4298, 
    3398, 
    3066, 
    2687, 
    6100, 
    3066, 
    6121, 
    3742, 
    1280, 
    4503, 
    4298, 
    3066, 
    6100, 
    4503, 
    3066, 
    5357, 
    6100, 
    2687, 
    4683, 
    4503, 
    6100, 
    781, 
    4980, 
    1357, 
    5450, 
    1615, 
    1027, 
    3130, 
    5450, 
    2767, 
    4980, 
    1615, 
    5450, 
    3130, 
    3454, 
    4649, 
    5875, 
    873, 
    1310, 
    1161, 
    5875, 
    3270, 
    3849, 
    873, 
    5875, 
    817, 
    4141, 
    1643, 
    5507, 
    873, 
    3849, 
    1615, 
    2039, 
    1385, 
    781, 
    873, 
    2039, 
    5503, 
    5066, 
    1626, 
    2695, 
    5503, 
    1145, 
    2695, 
    3071, 
    5503, 
    5332, 
    1041, 
    1804, 
    3080, 
    1214, 
    838, 
    982, 
    1479, 
    1214, 
    982, 
    666, 
    1479, 
    3872, 
    961, 
    850, 
    939, 
    3872, 
    1724, 
    1746, 
    961, 
    3872, 
    3565, 
    1914, 
    1196, 
    1291, 
    2456, 
    1192, 
    1291, 
    4796, 
    2456, 
    3565, 
    4543, 
    1746, 
    2322, 
    1338, 
    2224, 
    1196, 
    2322, 
    2224, 
    3220, 
    2452, 
    2750, 
    4982, 
    3220, 
    2870, 
    1817, 
    4982, 
    2870, 
    2913, 
    3255, 
    4982, 
    3985, 
    2452, 
    3220, 
    2452, 
    3985, 
    1011, 
    3985, 
    3220, 
    4982, 
    2322, 
    3985, 
    3255, 
    1785, 
    1011, 
    3985, 
    1338, 
    1666, 
    2224, 
    2039, 
    873, 
    5507, 
    1357, 
    873, 
    781, 
    1357, 
    1310, 
    873, 
    5450, 
    3130, 
    4827, 
    4408, 
    3409, 
    3080, 
    5986, 
    4408, 
    3080, 
    3066, 
    6179, 
    2687, 
    3066, 
    6374, 
    6179, 
    4192, 
    3706, 
    4408, 
    6179, 
    5933, 
    5799, 
    4408, 
    6179, 
    4192, 
    5986, 
    2687, 
    6179, 
    5645, 
    2704, 
    3706, 
    3961, 
    5645, 
    4192, 
    3961, 
    1628, 
    5645, 
    1628, 
    799, 
    5645, 
    2704, 
    609, 
    5005, 
    6392, 
    4683, 
    6100, 
    5357, 
    6392, 
    6100, 
    1310, 
    1357, 
    6392, 
    1453, 
    4406, 
    4605, 
    5357, 
    838, 
    6392, 
    6235, 
    4860, 
    949, 
    4605, 
    6235, 
    1104, 
    4605, 
    5933, 
    6235, 
    1453, 
    4605, 
    1104, 
    4406, 
    3961, 
    5799, 
    4860, 
    1737, 
    949, 
    4860, 
    3693, 
    1737, 
    1104, 
    6235, 
    949, 
    4605, 
    5799, 
    5933, 
    1280, 
    5626, 
    6121, 
    4649, 
    3454, 
    3742, 
    6060, 
    4649, 
    6121, 
    4503, 
    6060, 
    4298, 
    4503, 
    4827, 
    6060, 
    4503, 
    4683, 
    4827, 
    5626, 
    1422, 
    1737, 
    3398, 
    6524, 
    3693, 
    1280, 
    1422, 
    5626, 
    3693, 
    5626, 
    1737, 
    838, 
    1214, 
    5332, 
    5332, 
    1214, 
    1041, 
    1161, 
    5332, 
    1804, 
    3270, 
    838, 
    5332, 
    2113, 
    3482, 
    3821, 
    1200, 
    1917, 
    1007, 
    4796, 
    1914, 
    2456, 
    2116, 
    2420, 
    1507, 
    2116, 
    1011, 
    2420, 
    1196, 
    4543, 
    3565, 
    1785, 
    2322, 
    1196, 
    4543, 
    961, 
    1746, 
    1666, 
    5265, 
    2224, 
    5363, 
    3310, 
    1465, 
    2224, 
    5265, 
    4543, 
    1666, 
    3617, 
    5265, 
    850, 
    2735, 
    3872, 
    3310, 
    4604, 
    1465, 
    5767, 
    1368, 
    6370, 
    1804, 
    5767, 
    1161, 
    5439, 
    1368, 
    5767, 
    4604, 
    5439, 
    2695, 
    3062, 
    1368, 
    5439, 
    3310, 
    3062, 
    4604, 
    850, 
    5363, 
    1465, 
    1666, 
    2012, 
    3617, 
    1643, 
    1368, 
    3062, 
    4141, 
    5507, 
    1643, 
    5767, 
    6370, 
    1161, 
    5767, 
    1804, 
    3071, 
    1341, 
    2326, 
    879, 
    6152, 
    2594, 
    3039, 
    3371, 
    6152, 
    3039, 
    3371, 
    4347, 
    6152, 
    5424, 
    4115, 
    3848, 
    2271, 
    5424, 
    3039, 
    1267, 
    4115, 
    5424, 
    4136, 
    2326, 
    1341, 
    3575, 
    3672, 
    3371, 
    3269, 
    2326, 
    4136, 
    2043, 
    2326, 
    1789, 
    4347, 
    4136, 
    5068, 
    6152, 
    4347, 
    2594, 
    3371, 
    3672, 
    4347, 
    4754, 
    1746, 
    3872, 
    4115, 
    1267, 
    1969, 
    738, 
    5099, 
    1969, 
    3848, 
    3371, 
    5424, 
    5068, 
    1341, 
    2015, 
    3504, 
    5197, 
    3188, 
    4136, 
    1341, 
    5068, 
    5197, 
    4347, 
    5068, 
    3188, 
    5197, 
    5068, 
    3504, 
    2838, 
    5197, 
    3672, 
    3269, 
    4136, 
    2594, 
    1724, 
    3039, 
    3872, 
    2271, 
    1724, 
    2735, 
    1267, 
    2271, 
    3872, 
    2735, 
    2271, 
    850, 
    1465, 
    2735, 
    899, 
    1789, 
    5879, 
    3699, 
    738, 
    1882, 
    1088, 
    2160, 
    1037, 
    5616, 
    3059, 
    4771, 
    1922, 
    6440, 
    4483, 
    2457, 
    3059, 
    5616, 
    1037, 
    2160, 
    1573, 
    3472, 
    4603, 
    6507, 
    6191, 
    1085, 
    2158, 
    626, 
    2401, 
    313, 
    3790, 
    4338, 
    1154, 
    314, 
    3509, 
    784, 
    312, 
    2401, 
    626, 
    4338, 
    311, 
    1154, 
    3509, 
    973, 
    784, 
    5729, 
    3790, 
    3863, 
    2401, 
    5729, 
    3509, 
    4338, 
    3790, 
    5729, 
    312, 
    4338, 
    2401, 
    312, 
    311, 
    4338, 
    3863, 
    4257, 
    3749, 
    2401, 
    4338, 
    5729, 
    1154, 
    2199, 
    4257, 
    310, 
    1154, 
    311, 
    4700, 
    5025, 
    2007, 
    928, 
    1636, 
    2199, 
    928, 
    1639, 
    1636, 
    1157, 
    4666, 
    928, 
    2032, 
    4911, 
    2551, 
    1334, 
    2010, 
    4911, 
    1334, 
    1857, 
    2010, 
    4873, 
    1988, 
    1302, 
    809, 
    2007, 
    5025, 
    6017, 
    1332, 
    2949, 
    2544, 
    6017, 
    2949, 
    4700, 
    1332, 
    6017, 
    4873, 
    4700, 
    4528, 
    2007, 
    1332, 
    4700, 
    3289, 
    4682, 
    772, 
    4682, 
    4297, 
    1988, 
    4013, 
    2678, 
    2341, 
    1045, 
    4992, 
    5095, 
    3058, 
    2678, 
    4013, 
    1942, 
    3687, 
    691, 
    5637, 
    5010, 
    2678, 
    3391, 
    6297, 
    3058, 
    5472, 
    2893, 
    5637, 
    5095, 
    4013, 
    1806, 
    4451, 
    4242, 
    4992, 
    3391, 
    3058, 
    4242, 
    5095, 
    4242, 
    4013, 
    1045, 
    5095, 
    1806, 
    4992, 
    4242, 
    5095, 
    309, 
    4992, 
    1045, 
    1543, 
    4451, 
    4992, 
    2551, 
    2341, 
    1370, 
    2032, 
    2551, 
    1370, 
    814, 
    1639, 
    2604, 
    2604, 
    1806, 
    2341, 
    2551, 
    2604, 
    2341, 
    1639, 
    928, 
    5104, 
    5104, 
    928, 
    4666, 
    1045, 
    5104, 
    4666, 
    2604, 
    1639, 
    5104, 
    309, 
    624, 
    4992, 
    181, 
    180, 
    1087, 
    953, 
    1087, 
    179, 
    953, 
    179, 
    178, 
    4864, 
    953, 
    1225, 
    182, 
    2090, 
    1457, 
    1087, 
    953, 
    2090, 
    181, 
    1087, 
    182, 
    180, 
    179, 
    1087, 
    4570, 
    178, 
    177, 
    176, 
    4745, 
    177, 
    2731, 
    3102, 
    4570, 
    4745, 
    2731, 
    4570, 
    1701, 
    4745, 
    176, 
    1701, 
    5296, 
    4745, 
    4531, 
    3238, 
    1041, 
    4876, 
    3549, 
    4705, 
    797, 
    1626, 
    3549, 
    4864, 
    1225, 
    1323, 
    953, 
    178, 
    1225, 
    1457, 
    608, 
    182, 
    1323, 
    682, 
    5563, 
    183, 
    608, 
    1457, 
    2090, 
    182, 
    1087, 
    1673, 
    863, 
    1420, 
    695, 
    4251, 
    5955, 
    3191, 
    863, 
    1673, 
    175, 
    1136, 
    1701, 
    6596, 
    173, 
    1136, 
    175, 
    6596, 
    1136, 
    175, 
    174, 
    6596, 
    1119, 
    1232, 
    303, 
    858, 
    2477, 
    2800, 
    4923, 
    1707, 
    913, 
    2686, 
    5851, 
    913, 
    749, 
    1976, 
    4923, 
    2726, 
    4109, 
    1951, 
    4923, 
    6070, 
    1707, 
    3681, 
    1244, 
    2258, 
    5018, 
    1277, 
    2280, 
    1707, 
    6070, 
    2258, 
    1976, 
    1277, 
    3681, 
    2351, 
    1976, 
    749, 
    1389, 
    1277, 
    1976, 
    2351, 
    1389, 
    1976, 
    1819, 
    2351, 
    749, 
    1247, 
    2261, 
    2351, 
    3727, 
    916, 
    2065, 
    2041, 
    3727, 
    877, 
    2041, 
    3119, 
    3727, 
    2351, 
    2261, 
    1389, 
    5031, 
    1392, 
    2353, 
    1710, 
    5031, 
    2353, 
    2261, 
    1247, 
    6314, 
    3119, 
    2261, 
    1710, 
    3727, 
    3119, 
    1710, 
    1389, 
    2261, 
    3119, 
    1247, 
    5217, 
    6314, 
    4732, 
    1734, 
    947, 
    1244, 
    5018, 
    1951, 
    2280, 
    1734, 
    4732, 
    2041, 
    2280, 
    1277, 
    877, 
    1734, 
    2280, 
    5010, 
    2032, 
    1370, 
    5285, 
    4090, 
    3052, 
    4368, 
    5285, 
    2671, 
    3548, 
    4090, 
    5285, 
    3052, 
    2258, 
    1244, 
    4368, 
    5952, 
    5285, 
    4090, 
    2258, 
    3052, 
    2477, 
    858, 
    2032, 
    2116, 
    1507, 
    1511, 
    4493, 
    5125, 
    3116, 
    1011, 
    1914, 
    2420, 
    2320, 
    1111, 
    1334, 
    1007, 
    1783, 
    1200, 
    1007, 
    1597, 
    4824, 
    3482, 
    1507, 
    4796, 
    761, 
    3482, 
    1982, 
    2113, 
    1507, 
    3482, 
    1917, 
    2113, 
    1007, 
    2423, 
    1511, 
    1507, 
    1917, 
    2423, 
    2113, 
    4066, 
    3098, 
    2726, 
    5125, 
    2444, 
    4843, 
    1917, 
    3213, 
    2423, 
    3213, 
    3426, 
    2444, 
    2423, 
    3213, 
    2863, 
    1917, 
    1200, 
    5024, 
    4696, 
    1200, 
    2226, 
    1668, 
    5256, 
    2226, 
    4520, 
    5967, 
    5024, 
    2444, 
    3426, 
    3098, 
    5024, 
    1200, 
    4696, 
    4520, 
    5024, 
    4696, 
    3213, 
    1917, 
    5024, 
    2113, 
    2423, 
    1507, 
    2726, 
    1951, 
    709, 
    4066, 
    2726, 
    709, 
    1552, 
    4066, 
    709, 
    4843, 
    2444, 
    3098, 
    3996, 
    4843, 
    4066, 
    3996, 
    2750, 
    5125, 
    2863, 
    3213, 
    2444, 
    6234, 
    4109, 
    2726, 
    3098, 
    6234, 
    2726, 
    4323, 
    4109, 
    6234, 
    4109, 
    3052, 
    1244, 
    3098, 
    4323, 
    6234, 
    2671, 
    3052, 
    4109, 
    2863, 
    1511, 
    2423, 
    5305, 
    2750, 
    3996, 
    2116, 
    3116, 
    1011, 
    4493, 
    1511, 
    2863, 
    2444, 
    4493, 
    2863, 
    3116, 
    2116, 
    4493, 
    2452, 
    3116, 
    2750, 
    2116, 
    1511, 
    4493, 
    5305, 
    3996, 
    2144, 
    1060, 
    5305, 
    2144, 
    2870, 
    3220, 
    5305, 
    709, 
    4285, 
    5833, 
    4256, 
    1451, 
    3429, 
    709, 
    5833, 
    1552, 
    5833, 
    1216, 
    4256, 
    2456, 
    1746, 
    1192, 
    2320, 
    4824, 
    1111, 
    3821, 
    1597, 
    1007, 
    2113, 
    3821, 
    1007, 
    761, 
    1597, 
    3821, 
    5240, 
    2473, 
    1866, 
    761, 
    3235, 
    6209, 
    761, 
    1982, 
    3235, 
    4451, 
    3391, 
    4242, 
    691, 
    4451, 
    1543, 
    691, 
    3687, 
    4451, 
    2678, 
    1370, 
    2341, 
    4911, 
    2032, 
    858, 
    2546, 
    4911, 
    858, 
    2010, 
    2551, 
    4911, 
    2010, 
    814, 
    2551, 
    1806, 
    2604, 
    5104, 
    2551, 
    814, 
    2604, 
    814, 
    809, 
    1639, 
    4528, 
    2544, 
    772, 
    5164, 
    2010, 
    1857, 
    814, 
    5164, 
    2007, 
    814, 
    2010, 
    5164, 
    4646, 
    3413, 
    3086, 
    5240, 
    4646, 
    4465, 
    2180, 
    3413, 
    4646, 
    3413, 
    2544, 
    2949, 
    4465, 
    4646, 
    3086, 
    1607, 
    2544, 
    3413, 
    772, 
    2544, 
    1607, 
    1332, 
    1857, 
    2318, 
    1111, 
    4824, 
    1781, 
    4824, 
    1597, 
    1004, 
    1781, 
    4824, 
    1004, 
    1783, 
    1007, 
    4824, 
    1966, 
    735, 
    2125, 
    1265, 
    1966, 
    1028, 
    2408, 
    1896, 
    735, 
    1483, 
    2408, 
    1966, 
    1483, 
    3289, 
    4615, 
    6209, 
    3235, 
    5240, 
    1597, 
    6209, 
    1004, 
    1597, 
    761, 
    6209, 
    2383, 
    2473, 
    4135, 
    3344, 
    2383, 
    1443, 
    3648, 
    5243, 
    1443, 
    6079, 
    6398, 
    5182, 
    2079, 
    3648, 
    1443, 
    6398, 
    2158, 
    1166, 
    3009, 
    6191, 
    6079, 
    2622, 
    1085, 
    6191, 
    3648, 
    2838, 
    3504, 
    822, 
    1085, 
    2622, 
    3874, 
    3235, 
    1982, 
    1866, 
    2473, 
    2383, 
    5240, 
    1122, 
    4646, 
    1045, 
    4666, 
    309, 
    809, 
    1636, 
    1639, 
    2301, 
    2293, 
    1765, 
    936, 
    2301, 
    1765, 
    1311, 
    1758, 
    2301, 
    3509, 
    3863, 
    973, 
    2293, 
    1302, 
    1765, 
    3863, 
    3790, 
    4257, 
    1758, 
    3863, 
    3749, 
    1758, 
    973, 
    3863, 
    3749, 
    1302, 
    2293, 
    6706, 
    300, 
    1119, 
    301, 
    6706, 
    302, 
    301, 
    300, 
    6706, 
    300, 
    299, 
    1119, 
    3030, 
    299, 
    298, 
    6252, 
    2686, 
    2062, 
    6032, 
    5432, 
    4861, 
    2168, 
    2686, 
    5432, 
    4402, 
    4188, 
    3026, 
    913, 
    4402, 
    2062, 
    5817, 
    3548, 
    5669, 
    1707, 
    3823, 
    913, 
    5669, 
    3237, 
    5472, 
    6031, 
    4188, 
    5817, 
    1707, 
    2258, 
    4090, 
    5285, 
    3052, 
    2671, 
    3823, 
    4090, 
    3548, 
    3823, 
    1707, 
    4090, 
    2893, 
    5010, 
    5637, 
    3026, 
    1414, 
    2062, 
    913, 
    3823, 
    4402, 
    5819, 
    1119, 
    299, 
    1414, 
    5819, 
    299, 
    3358, 
    1119, 
    5819, 
    4188, 
    3955, 
    3358, 
    2062, 
    4402, 
    3026, 
    5817, 
    3823, 
    3548, 
    1232, 
    1119, 
    3358, 
    3026, 
    3358, 
    5819, 
    302, 
    1119, 
    303, 
    302, 
    6706, 
    1119, 
    5285, 
    3237, 
    3548, 
    5866, 
    4368, 
    2671, 
    4323, 
    5866, 
    2671, 
    4323, 
    4520, 
    5866, 
    5952, 
    3237, 
    5285, 
    4157, 
    5952, 
    4368, 
    4157, 
    2893, 
    5952, 
    5010, 
    2893, 
    2477, 
    2032, 
    5010, 
    2477, 
    2678, 
    3058, 
    5637, 
    3955, 
    1232, 
    3358, 
    4242, 
    3058, 
    4013, 
    3687, 
    3391, 
    4451, 
    1232, 
    3955, 
    1942, 
    5817, 
    4188, 
    4402, 
    3823, 
    5817, 
    4402, 
    6529, 
    5472, 
    6297, 
    3237, 
    5669, 
    3548, 
    6297, 
    3391, 
    5903, 
    6529, 
    6297, 
    5903, 
    5472, 
    5637, 
    6297, 
    2893, 
    5472, 
    3237, 
    5903, 
    3687, 
    3955, 
    6529, 
    5903, 
    6031, 
    5817, 
    6529, 
    6031, 
    5669, 
    5472, 
    6529, 
    3391, 
    3687, 
    5903, 
    1942, 
    3955, 
    3687, 
    3358, 
    3026, 
    4188, 
    6297, 
    5637, 
    3058, 
    307, 
    6658, 
    691, 
    304, 
    1232, 
    1942, 
    3026, 
    5819, 
    1414, 
    1543, 
    623, 
    691, 
    305, 
    6603, 
    306, 
    6658, 
    304, 
    1942, 
    6603, 
    6658, 
    307, 
    6603, 
    304, 
    6658, 
    306, 
    6603, 
    307, 
    305, 
    304, 
    6603, 
    6658, 
    1942, 
    691, 
    307, 
    691, 
    623, 
    308, 
    623, 
    1543, 
    1819, 
    6265, 
    1954, 
    2351, 
    1819, 
    1247, 
    1583, 
    2168, 
    6265, 
    5851, 
    2686, 
    1583, 
    749, 
    5851, 
    1583, 
    4923, 
    913, 
    5851, 
    2168, 
    5152, 
    6265, 
    4876, 
    5563, 
    682, 
    5563, 
    4864, 
    1323, 
    4531, 
    5775, 
    5911, 
    1457, 
    2090, 
    5027, 
    2090, 
    953, 
    4864, 
    1785, 
    1196, 
    1914, 
    5529, 
    1385, 
    3886, 
    4801, 
    5529, 
    3886, 
    2913, 
    2349, 
    5529, 
    1132, 
    2349, 
    1817, 
    4350, 
    1027, 
    1615, 
    1132, 
    4350, 
    2349, 
    1132, 
    1027, 
    4350, 
    5363, 
    4543, 
    5265, 
    2012, 
    1666, 
    1338, 
    3255, 
    4801, 
    1338, 
    817, 
    3617, 
    2012, 
    3617, 
    3062, 
    3310, 
    5265, 
    3617, 
    3310, 
    817, 
    1643, 
    3617, 
    5164, 
    1857, 
    1332, 
    2546, 
    1334, 
    4911, 
    1668, 
    2546, 
    858, 
    1668, 
    2226, 
    2546, 
    5164, 
    1332, 
    2007, 
    1111, 
    1857, 
    1334, 
    1111, 
    1781, 
    2318, 
    2546, 
    2226, 
    2320, 
    1857, 
    1111, 
    2318, 
    3030, 
    1414, 
    299, 
    6032, 
    4861, 
    3030, 
    296, 
    6032, 
    297, 
    296, 
    1097, 
    6032, 
    6252, 
    5432, 
    2686, 
    1414, 
    6252, 
    2062, 
    4861, 
    5432, 
    6252, 
    297, 
    6032, 
    3030, 
    1097, 
    2168, 
    5432, 
    6031, 
    3955, 
    4188, 
    5669, 
    6529, 
    5817, 
    5903, 
    3955, 
    6031, 
    1370, 
    2678, 
    5010, 
    2341, 
    1806, 
    4013, 
    624, 
    1543, 
    4992, 
    624, 
    308, 
    1543, 
    304, 
    303, 
    1232, 
    1555, 
    1097, 
    6667, 
    297, 
    3030, 
    298, 
    6032, 
    1097, 
    5432, 
    1555, 
    294, 
    293, 
    5599, 
    1687, 
    3382, 
    5152, 
    2168, 
    1097, 
    713, 
    5152, 
    1555, 
    6265, 
    1819, 
    1583, 
    713, 
    6265, 
    5152, 
    713, 
    1954, 
    6265, 
    4053, 
    3321, 
    5909, 
    1068, 
    4053, 
    280, 
    1068, 
    3630, 
    4053, 
    1964, 
    1187, 
    5710, 
    1612, 
    622, 
    769, 
    4923, 
    5851, 
    749, 
    1414, 
    4861, 
    6252, 
    2168, 
    1583, 
    2686, 
    1414, 
    3030, 
    4861, 
    1097, 
    1555, 
    5152, 
    6667, 
    1097, 
    296, 
    2686, 
    913, 
    2062, 
    1954, 
    1247, 
    1819, 
    3382, 
    5032, 
    713, 
    5032, 
    2045, 
    5217, 
    2226, 
    1200, 
    1783, 
    2320, 
    2226, 
    1783, 
    4824, 
    2320, 
    1783, 
    1334, 
    2546, 
    2320, 
    1951, 
    4109, 
    1244, 
    5256, 
    2800, 
    4157, 
    2800, 
    2477, 
    2893, 
    4157, 
    2800, 
    2893, 
    5866, 
    4520, 
    6145, 
    5256, 
    1668, 
    2800, 
    6145, 
    5256, 
    4157, 
    4696, 
    2226, 
    5256, 
    1668, 
    858, 
    2800, 
    5952, 
    2893, 
    3237, 
    6145, 
    4157, 
    4368, 
    5866, 
    6145, 
    4368, 
    4520, 
    4696, 
    6145, 
    5967, 
    4520, 
    4323, 
    3098, 
    5967, 
    4323, 
    3426, 
    5024, 
    5967, 
    4696, 
    5256, 
    6145, 
    6070, 
    1976, 
    3681, 
    2258, 
    6070, 
    3681, 
    4923, 
    1976, 
    6070, 
    4323, 
    2671, 
    4109, 
    3426, 
    5967, 
    3098, 
    3426, 
    3213, 
    5024, 
    6667, 
    295, 
    294, 
    1555, 
    6667, 
    294, 
    296, 
    295, 
    6667, 
    1823, 
    4111, 
    3844, 
    916, 
    1823, 
    1066, 
    2353, 
    1392, 
    4795, 
    1710, 
    2353, 
    1823, 
    1710, 
    2261, 
    5031, 
    5823, 
    2387, 
    881, 
    6223, 
    5962, 
    3925, 
    5962, 
    5710, 
    2387, 
    3653, 
    6223, 
    3925, 
    5049, 
    4905, 
    5962, 
    4194, 
    4148, 
    5789, 
    2690, 
    4194, 
    2784, 
    5900, 
    2662, 
    4905, 
    945, 
    1964, 
    2662, 
    4930, 
    682, 
    3431, 
    3102, 
    5069, 
    3431, 
    2797, 
    1088, 
    4757, 
    4757, 
    797, 
    682, 
    6440, 
    1516, 
    5616, 
    4483, 
    6440, 
    5616, 
    1064, 
    1516, 
    6440, 
    1037, 
    1626, 
    1088, 
    1145, 
    1037, 
    1573, 
    1366, 
    1882, 
    738, 
    1969, 
    1366, 
    738, 
    6112, 
    4806, 
    4698, 
    5668, 
    6112, 
    3848, 
    5668, 
    4959, 
    6112, 
    5099, 
    4959, 
    5668, 
    1969, 
    5099, 
    4115, 
    738, 
    4074, 
    5099, 
    4074, 
    3689, 
    4959, 
    4806, 
    4959, 
    3392, 
    1573, 
    4074, 
    738, 
    1573, 
    3957, 
    4074, 
    1516, 
    1699, 
    2457, 
    1267, 
    2735, 
    5859, 
    3062, 
    3617, 
    1643, 
    1969, 
    1267, 
    5859, 
    5363, 
    850, 
    961, 
    4543, 
    5363, 
    961, 
    5265, 
    3310, 
    5363, 
    1882, 
    4604, 
    2695, 
    3699, 
    1882, 
    1145, 
    1573, 
    3699, 
    1145, 
    1573, 
    738, 
    3699, 
    4604, 
    3062, 
    5439, 
    1366, 
    4604, 
    1882, 
    1366, 
    1465, 
    4604, 
    3270, 
    5875, 
    1310, 
    838, 
    3270, 
    1310, 
    6370, 
    1368, 
    1643, 
    5875, 
    6370, 
    3849, 
    5875, 
    1161, 
    6370, 
    5332, 
    1161, 
    3270, 
    5582, 
    3071, 
    1804, 
    1041, 
    5582, 
    1804, 
    3238, 
    5066, 
    5582, 
    3071, 
    5439, 
    5767, 
    3071, 
    2695, 
    5439, 
    1041, 
    3238, 
    5582, 
    5066, 
    5503, 
    3071, 
    1145, 
    1882, 
    2695, 
    6370, 
    1643, 
    3849, 
    5911, 
    4705, 
    4531, 
    1457, 
    5911, 
    5775, 
    5027, 
    5563, 
    5911, 
    5563, 
    4705, 
    5911, 
    4864, 
    5563, 
    5027, 
    4876, 
    4705, 
    5563, 
    797, 
    4876, 
    682, 
    797, 
    3549, 
    4876, 
    3549, 
    3238, 
    4705, 
    6707, 
    292, 
    291, 
    5599, 
    291, 
    1687, 
    1555, 
    5599, 
    3382, 
    6707, 
    291, 
    5599, 
    293, 
    6707, 
    5599, 
    293, 
    292, 
    6707, 
    279, 
    278, 
    6647, 
    267, 
    1189, 
    268, 
    269, 
    268, 
    1189, 
    6629, 
    273, 
    272, 
    6570, 
    6629, 
    272, 
    274, 
    273, 
    6629, 
    6570, 
    272, 
    6569, 
    274, 
    6629, 
    620, 
    620, 
    6629, 
    6570, 
    6569, 
    272, 
    271, 
    6569, 
    620, 
    6570, 
    2677, 
    6628, 
    271, 
    275, 
    620, 
    6569, 
    847, 
    1800, 
    2677, 
    1210, 
    277, 
    276, 
    1800, 
    1210, 
    276, 
    2677, 
    1800, 
    275, 
    6628, 
    2677, 
    275, 
    6569, 
    6628, 
    275, 
    6569, 
    271, 
    6628, 
    271, 
    3572, 
    2677, 
    5205, 
    6348, 
    2865, 
    271, 
    619, 
    3572, 
    1661, 
    619, 
    270, 
    2429, 
    2703, 
    3408, 
    270, 
    2221, 
    1661, 
    269, 
    1189, 
    2221, 
    2291, 
    1068, 
    6647, 
    1958, 
    3695, 
    719, 
    1006, 
    2592, 
    778, 
    5338, 
    3630, 
    2148, 
    1560, 
    5338, 
    2148, 
    5760, 
    6536, 
    5595, 
    5789, 
    4148, 
    3695, 
    3465, 
    5789, 
    3695, 
    3143, 
    2784, 
    5789, 
    6202, 
    4148, 
    5595, 
    5338, 
    6202, 
    6085, 
    3898, 
    4148, 
    6202, 
    2291, 
    2148, 
    1068, 
    1756, 
    1560, 
    2148, 
    1210, 
    4978, 
    2291, 
    6348, 
    5218, 
    5970, 
    2865, 
    6348, 
    5970, 
    5205, 
    5871, 
    6348, 
    3962, 
    1731, 
    945, 
    5338, 
    6085, 
    3630, 
    3465, 
    1958, 
    1251, 
    4629, 
    3465, 
    1251, 
    870, 
    4629, 
    1251, 
    3070, 
    2694, 
    4802, 
    3695, 
    3898, 
    719, 
    3143, 
    5789, 
    3465, 
    5789, 
    2784, 
    4194, 
    5973, 
    5049, 
    5183, 
    3321, 
    3630, 
    6085, 
    5595, 
    5900, 
    5760, 
    6536, 
    6202, 
    5595, 
    3321, 
    6085, 
    5973, 
    5338, 
    3898, 
    6202, 
    4148, 
    4194, 
    5595, 
    3695, 
    4148, 
    3898, 
    5900, 
    3962, 
    2662, 
    3695, 
    1958, 
    3465, 
    2429, 
    1319, 
    1520, 
    2703, 
    2429, 
    1520, 
    2120, 
    4845, 
    6196, 
    4069, 
    2221, 
    3079, 
    3408, 
    4288, 
    3079, 
    2447, 
    1661, 
    4069, 
    1924, 
    1206, 
    2429, 
    266, 
    265, 
    6701, 
    6662, 
    213, 
    212, 
    211, 
    6662, 
    212, 
    211, 
    758, 
    6662, 
    6662, 
    758, 
    213, 
    6651, 
    220, 
    6593, 
    6703, 
    219, 
    218, 
    6593, 
    6703, 
    218, 
    220, 
    219, 
    6703, 
    218, 
    6592, 
    6593, 
    6593, 
    220, 
    6703, 
    223, 
    6593, 
    6592, 
    6651, 
    221, 
    220, 
    222, 
    6651, 
    6593, 
    222, 
    221, 
    6651, 
    718, 
    218, 
    614, 
    217, 
    216, 
    1559, 
    1559, 
    216, 
    1168, 
    614, 
    1559, 
    718, 
    614, 
    217, 
    1559, 
    2209, 
    1648, 
    1168, 
    6593, 
    223, 
    222, 
    1957, 
    6592, 
    218, 
    1957, 
    223, 
    6592, 
    718, 
    1957, 
    218, 
    718, 
    1897, 
    1957, 
    215, 
    2209, 
    216, 
    1252, 
    5578, 
    1854, 
    5015, 
    4660, 
    720, 
    1854, 
    5578, 
    720, 
    6033, 
    4838, 
    4660, 
    4226, 
    6033, 
    5015, 
    4226, 
    2428, 
    6033, 
    1559, 
    1168, 
    1897, 
    2209, 
    214, 
    1648, 
    216, 
    2209, 
    1168, 
    215, 
    214, 
    2209, 
    1648, 
    758, 
    1594, 
    6612, 
    245, 
    1160, 
    246, 
    6612, 
    247, 
    246, 
    245, 
    6612, 
    243, 
    242, 
    1887, 
    242, 
    241, 
    1887, 
    6692, 
    238, 
    237, 
    6708, 
    237, 
    785, 
    6692, 
    6708, 
    240, 
    6692, 
    237, 
    6708, 
    239, 
    6692, 
    240, 
    239, 
    238, 
    6692, 
    236, 
    235, 
    6675, 
    6675, 
    235, 
    2397, 
    237, 
    6675, 
    785, 
    237, 
    236, 
    6675, 
    2397, 
    234, 
    233, 
    1995, 
    233, 
    232, 
    2566, 
    1150, 
    1995, 
    232, 
    2566, 
    1995, 
    1160, 
    244, 
    2566, 
    6708, 
    785, 
    240, 
    2397, 
    233, 
    1995, 
    785, 
    2397, 
    1995, 
    235, 
    234, 
    2397, 
    1150, 
    240, 
    785, 
    2397, 
    785, 
    6675, 
    1768, 
    2566, 
    232, 
    1150, 
    785, 
    1995, 
    1887, 
    1150, 
    244, 
    243, 
    1887, 
    244, 
    241, 
    1150, 
    1887, 
    241, 
    240, 
    1150, 
    1160, 
    987, 
    6612, 
    1150, 
    2566, 
    244, 
    1160, 
    2566, 
    1768, 
    987, 
    2239, 
    1016, 
    244, 
    1160, 
    245, 
    2239, 
    1688, 
    5259, 
    1016, 
    2239, 
    675, 
    1768, 
    232, 
    2239, 
    1160, 
    1768, 
    987, 
    232, 
    1688, 
    2239, 
    6594, 
    229, 
    1688, 
    230, 
    6594, 
    231, 
    230, 
    229, 
    6594, 
    1688, 
    231, 
    6594, 
    882, 
    5355, 
    229, 
    2239, 
    987, 
    1768, 
    231, 
    1688, 
    232, 
    6685, 
    616, 
    6676, 
    6685, 
    226, 
    616, 
    227, 
    6685, 
    6676, 
    227, 
    226, 
    6685, 
    882, 
    6676, 
    225, 
    6676, 
    228, 
    227, 
    225, 
    6676, 
    616, 
    882, 
    228, 
    6676, 
    2127, 
    225, 
    1923, 
    5259, 
    5355, 
    2127, 
    229, 
    228, 
    882, 
    6681, 
    224, 
    615, 
    6680, 
    6681, 
    615, 
    225, 
    224, 
    6681, 
    6680, 
    615, 
    223, 
    1923, 
    6680, 
    223, 
    225, 
    6681, 
    6680, 
    1897, 
    4660, 
    5196, 
    1559, 
    1897, 
    718, 
    4984, 
    824, 
    4660, 
    1897, 
    4984, 
    4660, 
    1168, 
    1648, 
    4984, 
    6612, 
    987, 
    247, 
    225, 
    6680, 
    1923, 
    4226, 
    5015, 
    5578, 
    1517, 
    4226, 
    3735, 
    6033, 
    1923, 
    4838, 
    213, 
    758, 
    214, 
    5912, 
    827, 
    1052, 
    5259, 
    675, 
    2239, 
    5355, 
    5259, 
    1688, 
    229, 
    5355, 
    1688, 
    882, 
    2127, 
    5355, 
    1517, 
    675, 
    5259, 
    2127, 
    2428, 
    5259, 
    225, 
    2127, 
    882, 
    2428, 
    1517, 
    5259, 
    1923, 
    2428, 
    2127, 
    4838, 
    5196, 
    4660, 
    5196, 
    4838, 
    1923, 
    1957, 
    5196, 
    223, 
    1957, 
    1897, 
    5196, 
    4660, 
    824, 
    720, 
    6033, 
    4660, 
    5015, 
    2428, 
    1923, 
    6033, 
    1923, 
    223, 
    5196, 
    1897, 
    1168, 
    4984, 
    1252, 
    1428, 
    2327, 
    247, 
    1016, 
    922, 
    247, 
    987, 
    1016, 
    2285, 
    1288, 
    2253, 
    2588, 
    2285, 
    1743, 
    3626, 
    1288, 
    2285, 
    1648, 
    1594, 
    824, 
    4984, 
    1648, 
    824, 
    214, 
    758, 
    1648, 
    758, 
    1288, 
    1594, 
    210, 
    904, 
    211, 
    1171, 
    700, 
    957, 
    1743, 
    1238, 
    1171, 
    4122, 
    2531, 
    2938, 
    2981, 
    4122, 
    3858, 
    6150, 
    2531, 
    4122, 
    957, 
    6150, 
    4122, 
    957, 
    700, 
    6150, 
    3626, 
    1594, 
    1288, 
    3626, 
    2174, 
    1594, 
    2588, 
    3626, 
    2285, 
    2588, 
    2981, 
    5593, 
    720, 
    824, 
    2174, 
    4295, 
    2850, 
    1591, 
    1330, 
    4295, 
    1591, 
    2712, 
    1171, 
    4295, 
    617, 
    829, 
    4669, 
    5902, 
    2938, 
    6255, 
    6217, 
    6399, 
    5902, 
    5707, 
    1252, 
    1854, 
    1428, 
    5707, 
    3279, 
    1428, 
    1252, 
    5707, 
    617, 
    833, 
    829, 
    6217, 
    922, 
    1715, 
    833, 
    5146, 
    3381, 
    248, 
    922, 
    5146, 
    6630, 
    261, 
    2244, 
    262, 
    6630, 
    263, 
    262, 
    261, 
    6630, 
    261, 
    1487, 
    2244, 
    737, 
    257, 
    256, 
    737, 
    258, 
    257, 
    5206, 
    1495, 
    737, 
    5206, 
    2414, 
    1495, 
    255, 
    5206, 
    256, 
    4580, 
    2414, 
    5206, 
    1906, 
    839, 
    2414, 
    4580, 
    1906, 
    2414, 
    254, 
    4580, 
    255, 
    254, 
    2153, 
    4580, 
    259, 
    258, 
    737, 
    251, 
    1182, 
    252, 
    1182, 
    2153, 
    252, 
    250, 
    1831, 
    251, 
    2153, 
    254, 
    253, 
    1297, 
    1906, 
    1182, 
    839, 
    1752, 
    3879, 
    2153, 
    1182, 
    1906, 
    4580, 
    2153, 
    1906, 
    253, 
    252, 
    2153, 
    5206, 
    255, 
    4580, 
    260, 
    618, 
    4267, 
    5943, 
    4267, 
    618, 
    1495, 
    5943, 
    259, 
    1495, 
    3879, 
    5943, 
    1495, 
    259, 
    737, 
    256, 
    5206, 
    737, 
    3879, 
    1752, 
    968, 
    2414, 
    3879, 
    1495, 
    2414, 
    839, 
    3879, 
    1831, 
    1297, 
    1182, 
    4669, 
    1831, 
    250, 
    1651, 
    1176, 
    2613, 
    5688, 
    1176, 
    1173, 
    1831, 
    2613, 
    1297, 
    1831, 
    4669, 
    2613, 
    4669, 
    1651, 
    2613, 
    3001, 
    1879, 
    1142, 
    4086, 
    3337, 
    3001, 
    2329, 
    6114, 
    1142, 
    6114, 
    1622, 
    5609, 
    5704, 
    6002, 
    4995, 
    3028, 
    2642, 
    3337, 
    3913, 
    3028, 
    3544, 
    829, 
    3360, 
    1651, 
    829, 
    833, 
    3381, 
    3360, 
    829, 
    3381, 
    3028, 
    3360, 
    5991, 
    5943, 
    3879, 
    968, 
    4267, 
    968, 
    261, 
    259, 
    5943, 
    618, 
    5943, 
    968, 
    4267, 
    1398, 
    2049, 
    839, 
    891, 
    968, 
    1752, 
    891, 
    1487, 
    968, 
    5688, 
    1173, 
    1398, 
    1487, 
    891, 
    1490, 
    2720, 
    1487, 
    1490, 
    4952, 
    2720, 
    1490, 
    1900, 
    4952, 
    1490, 
    2590, 
    793, 
    4952, 
    1676, 
    1319, 
    2720, 
    2244, 
    263, 
    6630, 
    991, 
    2244, 
    1487, 
    991, 
    264, 
    2244, 
    2720, 
    991, 
    1487, 
    1019, 
    2120, 
    793, 
    1206, 
    991, 
    1319, 
    1924, 
    1189, 
    267, 
    1319, 
    2429, 
    1206, 
    4997, 
    5941, 
    6201, 
    6196, 
    6201, 
    6292, 
    2447, 
    5479, 
    2865, 
    2447, 
    4069, 
    5479, 
    4069, 
    3079, 
    4288, 
    1189, 
    3408, 
    3079, 
    1924, 
    2429, 
    3408, 
    1676, 
    1520, 
    1319, 
    991, 
    2720, 
    1319, 
    793, 
    2120, 
    1676, 
    3408, 
    2703, 
    4288, 
    6201, 
    4845, 
    4997, 
    1520, 
    6196, 
    2703, 
    1520, 
    2120, 
    6196, 
    5218, 
    4978, 
    1800, 
    5970, 
    5218, 
    847, 
    2447, 
    5970, 
    847, 
    2447, 
    2865, 
    5970, 
    6348, 
    5871, 
    4978, 
    3216, 
    5205, 
    2865, 
    6348, 
    4978, 
    5218, 
    2511, 
    5871, 
    5205, 
    2511, 
    6008, 
    5871, 
    719, 
    1560, 
    6008, 
    2922, 
    719, 
    6008, 
    1676, 
    2120, 
    1520, 
    1958, 
    2922, 
    6497, 
    6497, 
    6102, 
    3807, 
    1251, 
    6497, 
    3807, 
    1251, 
    1958, 
    6497, 
    4871, 
    5253, 
    5918, 
    5479, 
    6510, 
    2865, 
    5613, 
    6149, 
    2329, 
    6701, 
    267, 
    266, 
    1924, 
    6701, 
    265, 
    1924, 
    267, 
    6701, 
    264, 
    263, 
    2244, 
    261, 
    260, 
    4267, 
    2981, 
    3858, 
    5665, 
    5146, 
    833, 
    248, 
    6217, 
    3047, 
    3381, 
    922, 
    6217, 
    5146, 
    6399, 
    1428, 
    3279, 
    1715, 
    6399, 
    6217, 
    1715, 
    1428, 
    6399, 
    5991, 
    3360, 
    3381, 
    3047, 
    5991, 
    3381, 
    3047, 
    2665, 
    6493, 
    5146, 
    6217, 
    3381, 
    6493, 
    2642, 
    3028, 
    2665, 
    6002, 
    6493, 
    2665, 
    4995, 
    6002, 
    1715, 
    1016, 
    2327, 
    6493, 
    6002, 
    2642, 
    5991, 
    6493, 
    3028, 
    5991, 
    3047, 
    6493, 
    5902, 
    2665, 
    3047, 
    6217, 
    5902, 
    3047, 
    3279, 
    2938, 
    5902, 
    2531, 
    1461, 
    4995, 
    922, 
    1016, 
    1715, 
    5475, 
    3658, 
    4579, 
    1633, 
    5475, 
    4584, 
    3356, 
    3658, 
    5475, 
    1424, 
    3356, 
    5475, 
    5965, 
    4171, 
    1345, 
    827, 
    5965, 
    1052, 
    827, 
    4386, 
    5965, 
    5965, 
    4579, 
    4171, 
    6048, 
    4386, 
    827, 
    1548, 
    6048, 
    827, 
    1548, 
    5293, 
    6048, 
    4584, 
    5475, 
    4579, 
    6015, 
    2725, 
    921, 
    4871, 
    6015, 
    5021, 
    5023, 
    2725, 
    6015, 
    4699, 
    6503, 
    4871, 
    3658, 
    3356, 
    5023, 
    2725, 
    5023, 
    3356, 
    5253, 
    4871, 
    5021, 
    3216, 
    5807, 
    3528, 
    5918, 
    5445, 
    5613, 
    5253, 
    5847, 
    5140, 
    4845, 
    1019, 
    5445, 
    6195, 
    4699, 
    4527, 
    4171, 
    6195, 
    4527, 
    4171, 
    3931, 
    6195, 
    5021, 
    2400, 
    3807, 
    5023, 
    6015, 
    4871, 
    6015, 
    1714, 
    5021, 
    2329, 
    1142, 
    1345, 
    793, 
    1622, 
    1019, 
    5337, 
    2590, 
    2983, 
    5820, 
    5337, 
    2983, 
    3544, 
    3337, 
    5337, 
    5609, 
    3337, 
    4086, 
    1173, 
    5820, 
    2983, 
    1176, 
    1651, 
    3913, 
    2642, 
    3001, 
    3337, 
    6149, 
    1622, 
    1378, 
    793, 
    2720, 
    4952, 
    5902, 
    6399, 
    3279, 
    6255, 
    2531, 
    4995, 
    5902, 
    6255, 
    2665, 
    2938, 
    2531, 
    6255, 
    5665, 
    1854, 
    2981, 
    3279, 
    5707, 
    3858, 
    5707, 
    1854, 
    5665, 
    4122, 
    2588, 
    957, 
    4122, 
    2981, 
    2588, 
    3279, 
    3858, 
    2938, 
    3858, 
    5707, 
    5665, 
    1854, 
    720, 
    5593, 
    5704, 
    1879, 
    3001, 
    6255, 
    4995, 
    2665, 
    1461, 
    827, 
    5912, 
    4669, 
    829, 
    1651, 
    249, 
    4669, 
    250, 
    249, 
    617, 
    4669, 
    617, 
    248, 
    833, 
    1807, 
    209, 
    208, 
    5300, 
    3928, 
    1704, 
    1948, 
    5300, 
    910, 
    1002, 
    3928, 
    5300, 
    3928, 
    904, 
    210, 
    910, 
    5300, 
    1704, 
    1002, 
    904, 
    3928, 
    2240, 
    692, 
    1689, 
    2640, 
    2600, 
    1943, 
    2247, 
    5235, 
    1233, 
    2365, 
    1411, 
    3328, 
    3203, 
    5277, 
    910, 
    1233, 
    2640, 
    1943, 
    5277, 
    2059, 
    910, 
    2775, 
    5277, 
    3203, 
    3328, 
    2059, 
    5277, 
    756, 
    5300, 
    1948, 
    4295, 
    1330, 
    2712, 
    1948, 
    1591, 
    756, 
    706, 
    1330, 
    1591, 
    3928, 
    210, 
    209, 
    1807, 
    208, 
    207, 
    5993, 
    2775, 
    3203, 
    4218, 
    209, 
    1807, 
    4280, 
    4218, 
    1807, 
    1046, 
    4280, 
    1807, 
    6218, 
    3203, 
    910, 
    4280, 
    6218, 
    4218, 
    5993, 
    3203, 
    6218, 
    4059, 
    5993, 
    4280, 
    4059, 
    1544, 
    5993, 
    1704, 
    209, 
    4218, 
    922, 
    248, 
    247, 
    4108, 
    2327, 
    1016, 
    675, 
    4108, 
    1016, 
    675, 
    1517, 
    4108, 
    4226, 
    1517, 
    2428, 
    2327, 
    3735, 
    1252, 
    2327, 
    4108, 
    3735, 
    1715, 
    2327, 
    1428, 
    4108, 
    1517, 
    3735, 
    2588, 
    1743, 
    957, 
    4122, 
    2938, 
    3858, 
    5593, 
    2174, 
    3626, 
    2588, 
    5593, 
    3626, 
    2981, 
    1854, 
    5593, 
    5578, 
    5015, 
    720, 
    3735, 
    5578, 
    1252, 
    3735, 
    4226, 
    5578, 
    720, 
    2174, 
    5593, 
    4920, 
    5193, 
    5293, 
    1461, 
    1548, 
    827, 
    1461, 
    2531, 
    6150, 
    1548, 
    6150, 
    700, 
    1345, 
    1879, 
    1052, 
    1461, 
    6150, 
    1548, 
    2174, 
    824, 
    1594, 
    5204, 
    895, 
    2052, 
    2717, 
    3161, 
    1094, 
    2717, 
    1696, 
    3161, 
    1844, 
    2717, 
    1094, 
    2247, 
    1936, 
    677, 
    2717, 
    5235, 
    1696, 
    895, 
    3161, 
    1696, 
    1844, 
    2365, 
    5113, 
    1233, 
    1936, 
    2247, 
    6216, 
    2803, 
    3522, 
    2666, 
    6304, 
    6029, 
    2440, 
    2803, 
    6216, 
    2725, 
    2068, 
    921, 
    6029, 
    1815, 
    2666, 
    6304, 
    6216, 
    6029, 
    3048, 
    6304, 
    2666, 
    2440, 
    6216, 
    6304, 
    3522, 
    1424, 
    6029, 
    1105, 
    2142, 
    806, 
    6029, 
    1424, 
    1815, 
    5188, 
    3522, 
    2803, 
    2068, 
    1424, 
    3522, 
    3158, 
    2803, 
    2440, 
    1973, 
    3965, 
    746, 
    3965, 
    4913, 
    3158, 
    1633, 
    1815, 
    1424, 
    3048, 
    1094, 
    2165, 
    2440, 
    6304, 
    2165, 
    2666, 
    1057, 
    4612, 
    5204, 
    3161, 
    895, 
    2165, 
    1094, 
    3161, 
    5204, 
    2165, 
    3161, 
    1402, 
    5204, 
    2052, 
    1580, 
    2165, 
    5204, 
    2666, 
    1815, 
    1057, 
    2142, 
    4612, 
    1057, 
    6029, 
    6216, 
    3522, 
    1580, 
    2440, 
    2165, 
    1580, 
    746, 
    3158, 
    2571, 
    1550, 
    3635, 
    1844, 
    2571, 
    2365, 
    2142, 
    1550, 
    2571, 
    806, 
    2142, 
    1057, 
    1105, 
    1550, 
    2142, 
    1943, 
    2600, 
    692, 
    5113, 
    2717, 
    1844, 
    3328, 
    5113, 
    2365, 
    2640, 
    1233, 
    5235, 
    706, 
    1948, 
    2059, 
    1535, 
    677, 
    2919, 
    2291, 
    278, 
    1210, 
    1800, 
    4978, 
    1210, 
    1756, 
    2148, 
    2291, 
    968, 
    1487, 
    261, 
    2720, 
    793, 
    1676, 
    1752, 
    2049, 
    891, 
    1900, 
    2983, 
    4952, 
    2049, 
    1398, 
    1900, 
    891, 
    2049, 
    1900, 
    1752, 
    839, 
    2049, 
    1622, 
    2590, 
    5609, 
    1831, 
    1182, 
    251, 
    5688, 
    1297, 
    2613, 
    1176, 
    5688, 
    2613, 
    1398, 
    1297, 
    5688, 
    1900, 
    1398, 
    1173, 
    2983, 
    1900, 
    1173, 
    5820, 
    3544, 
    5337, 
    1176, 
    5820, 
    1173, 
    1176, 
    3544, 
    5820, 
    2590, 
    4952, 
    2983, 
    3544, 
    3028, 
    3337, 
    1622, 
    793, 
    2590, 
    1490, 
    891, 
    1900, 
    839, 
    1297, 
    1398, 
    839, 
    1906, 
    1297, 
    3913, 
    3360, 
    3028, 
    1176, 
    3913, 
    3544, 
    1651, 
    3360, 
    3913, 
    5293, 
    2712, 
    4920, 
    6334, 
    6048, 
    5293, 
    4584, 
    6334, 
    5193, 
    4386, 
    6048, 
    6334, 
    700, 
    1171, 
    5293, 
    6299, 
    2690, 
    2784, 
    4956, 
    6299, 
    2784, 
    4197, 
    2277, 
    6299, 
    847, 
    1661, 
    2447, 
    2400, 
    1714, 
    870, 
    3216, 
    2511, 
    5205, 
    6497, 
    2922, 
    6102, 
    1958, 
    719, 
    2922, 
    4527, 
    2329, 
    1345, 
    3658, 
    5023, 
    6503, 
    5847, 
    5941, 
    5140, 
    2865, 
    6510, 
    3216, 
    6292, 
    4288, 
    2703, 
    6196, 
    6292, 
    2703, 
    6554, 
    5941, 
    5807, 
    2725, 
    3356, 
    2068, 
    806, 
    1633, 
    4584, 
    806, 
    1057, 
    1633, 
    3048, 
    2165, 
    6304, 
    2068, 
    3356, 
    1424, 
    1633, 
    1057, 
    1815, 
    1206, 
    264, 
    991, 
    1206, 
    1924, 
    265, 
    6102, 
    2511, 
    3216, 
    3807, 
    6102, 
    3528, 
    2922, 
    2511, 
    6102, 
    2221, 
    4069, 
    1661, 
    6102, 
    3216, 
    3528, 
    2221, 
    270, 
    269, 
    5479, 
    4069, 
    4288, 
    1189, 
    3079, 
    2221, 
    1189, 
    1924, 
    3408, 
    3572, 
    619, 
    1661, 
    847, 
    3572, 
    1661, 
    847, 
    2677, 
    3572, 
    264, 
    1206, 
    265, 
    1948, 
    706, 
    1591, 
    1002, 
    5300, 
    756, 
    2059, 
    1411, 
    706, 
    910, 
    2059, 
    1948, 
    2775, 
    1544, 
    692, 
    3328, 
    5277, 
    2600, 
    6218, 
    1704, 
    4218, 
    2600, 
    5277, 
    2775, 
    910, 
    1704, 
    6218, 
    1006, 
    3794, 
    281, 
    6653, 
    284, 
    621, 
    283, 
    1569, 
    621, 
    1569, 
    286, 
    285, 
    6653, 
    1569, 
    285, 
    284, 
    6653, 
    285, 
    621, 
    1569, 
    6653, 
    6585, 
    287, 
    1569, 
    283, 
    6585, 
    1569, 
    283, 
    3794, 
    6585, 
    287, 
    286, 
    1569, 
    769, 
    6585, 
    3794, 
    3794, 
    283, 
    282, 
    281, 
    3794, 
    282, 
    1006, 
    769, 
    3794, 
    769, 
    778, 
    1612, 
    287, 
    769, 
    622, 
    1006, 
    778, 
    769, 
    287, 
    6585, 
    769, 
    281, 
    280, 
    4053, 
    281, 
    5909, 
    1006, 
    6647, 
    1068, 
    280, 
    279, 
    6647, 
    280, 
    278, 
    2291, 
    6647, 
    5909, 
    2592, 
    1006, 
    4053, 
    5909, 
    281, 
    3321, 
    2592, 
    5909, 
    3630, 
    3321, 
    4053, 
    2148, 
    3630, 
    1068, 
    5338, 
    1560, 
    3898, 
    3898, 
    1560, 
    719, 
    290, 
    289, 
    1129, 
    1129, 
    289, 
    288, 
    5281, 
    845, 
    1731, 
    5341, 
    2147, 
    1066, 
    4460, 
    4250, 
    5341, 
    1835, 
    4460, 
    1081, 
    5736, 
    1798, 
    2984, 
    1835, 
    5736, 
    4460, 
    1835, 
    2358, 
    5736, 
    5114, 
    5736, 
    2984, 
    3844, 
    845, 
    2026, 
    5341, 
    3844, 
    2026, 
    4460, 
    5341, 
    2026, 
    4250, 
    2147, 
    5341, 
    1066, 
    1823, 
    3844, 
    5341, 
    1066, 
    3844, 
    1081, 
    4460, 
    2026, 
    1558, 
    1418, 
    2147, 
    1849, 
    2370, 
    717, 
    1418, 
    2065, 
    2147, 
    916, 
    1710, 
    1823, 
    2147, 
    2065, 
    1066, 
    717, 
    2370, 
    1558, 
    1956, 
    1849, 
    717, 
    6088, 
    670, 
    1451, 
    1100, 
    2899, 
    1849, 
    3984, 
    3427, 
    3718, 
    752, 
    5246, 
    1586, 
    3130, 
    2767, 
    4896, 
    5840, 
    2899, 
    2483, 
    6088, 
    5840, 
    2483, 
    670, 
    6088, 
    2483, 
    1216, 
    2792, 
    6088, 
    6363, 
    1849, 
    2899, 
    3471, 
    6363, 
    5840, 
    3471, 
    2370, 
    6363, 
    1100, 
    2171, 
    3718, 
    6251, 
    947, 
    1683, 
    2041, 
    877, 
    2280, 
    3119, 
    2041, 
    1389, 
    1710, 
    916, 
    3727, 
    1734, 
    877, 
    1683, 
    2045, 
    881, 
    1187, 
    1392, 
    2045, 
    1187, 
    5217, 
    1247, 
    1954, 
    1392, 
    5217, 
    2045, 
    6314, 
    5031, 
    2261, 
    1392, 
    6314, 
    5217, 
    1392, 
    5031, 
    6314, 
    1392, 
    1187, 
    1964, 
    4111, 
    1823, 
    2353, 
    5217, 
    1954, 
    5032, 
    2041, 
    1277, 
    1389, 
    749, 
    1583, 
    1819, 
    3382, 
    1687, 
    881, 
    1555, 
    3382, 
    713, 
    1555, 
    293, 
    5599, 
    1612, 
    288, 
    622, 
    6223, 
    5049, 
    5962, 
    1612, 
    6223, 
    3653, 
    5183, 
    5049, 
    6223, 
    2592, 
    5183, 
    778, 
    5973, 
    5760, 
    5049, 
    2592, 
    5973, 
    5183, 
    2592, 
    3321, 
    5973, 
    3653, 
    288, 
    1612, 
    5823, 
    1129, 
    3925, 
    2387, 
    5823, 
    3925, 
    1687, 
    291, 
    5823, 
    5032, 
    3382, 
    881, 
    2045, 
    5032, 
    881, 
    1954, 
    713, 
    5032, 
    291, 
    1129, 
    5823, 
    291, 
    290, 
    1129, 
    1535, 
    895, 
    1696, 
    3744, 
    1081, 
    1274, 
    2358, 
    1835, 
    3744, 
    3478, 
    2358, 
    3744, 
    1402, 
    1798, 
    2358, 
    4460, 
    5736, 
    5114, 
    5757, 
    5225, 
    2593, 
    2129, 
    5322, 
    1033, 
    2129, 
    4330, 
    5322, 
    1558, 
    2147, 
    4250, 
    2129, 
    895, 
    1535, 
    1402, 
    2052, 
    1033, 
    1402, 
    3478, 
    5204, 
    1798, 
    1402, 
    1033, 
    3478, 
    1580, 
    5204, 
    2358, 
    3478, 
    1402, 
    746, 
    1580, 
    3478, 
    731, 
    945, 
    1731, 
    2712, 
    5293, 
    1171, 
    1238, 
    4295, 
    1171, 
    5193, 
    806, 
    4584, 
    1330, 
    4920, 
    2712, 
    1105, 
    806, 
    5193, 
    1550, 
    1105, 
    1330, 
    3635, 
    1550, 
    706, 
    1411, 
    3635, 
    706, 
    1411, 
    2365, 
    3635, 
    4612, 
    1094, 
    3048, 
    3635, 
    2365, 
    2571, 
    5235, 
    5113, 
    2640, 
    1696, 
    5235, 
    2247, 
    2717, 
    5113, 
    5235, 
    1094, 
    4612, 
    1844, 
    3328, 
    2600, 
    2640, 
    5113, 
    3328, 
    2640, 
    1411, 
    2059, 
    3328, 
    6334, 
    4584, 
    4386, 
    6334, 
    5293, 
    5193, 
    4920, 
    1105, 
    5193, 
    3522, 
    5188, 
    2068, 
    1580, 
    3158, 
    2440, 
    6327, 
    3070, 
    870, 
    921, 
    6327, 
    1714, 
    5188, 
    4913, 
    6327, 
    3158, 
    4913, 
    2803, 
    2694, 
    3070, 
    4913, 
    3962, 
    945, 
    2662, 
    6299, 
    1731, 
    2690, 
    4197, 
    1274, 
    2277, 
    5438, 
    2694, 
    3965, 
    1973, 
    5438, 
    3965, 
    4197, 
    4956, 
    5438, 
    1731, 
    6299, 
    2277, 
    4956, 
    4802, 
    2694, 
    6299, 
    4956, 
    4197, 
    2784, 
    3143, 
    4956, 
    3962, 
    4194, 
    2690, 
    1731, 
    3962, 
    2690, 
    5900, 
    4905, 
    5760, 
    4194, 
    5900, 
    5595, 
    4194, 
    3962, 
    5900, 
    4802, 
    3465, 
    4629, 
    5188, 
    6327, 
    921, 
    1274, 
    1081, 
    5281, 
    5281, 
    1081, 
    2026, 
    845, 
    5281, 
    2026, 
    2277, 
    1274, 
    5281, 
    4845, 
    2120, 
    1019, 
    5445, 
    4997, 
    4845, 
    6149, 
    5613, 
    5445, 
    1622, 
    6149, 
    1019, 
    1378, 
    2329, 
    6149, 
    5918, 
    4699, 
    4871, 
    4997, 
    5918, 
    5140, 
    5613, 
    4699, 
    5918, 
    6510, 
    5807, 
    3216, 
    6292, 
    6510, 
    5479, 
    6554, 
    6201, 
    5941, 
    6292, 
    6554, 
    6510, 
    6292, 
    6201, 
    6554, 
    6510, 
    6554, 
    5807, 
    4288, 
    6292, 
    5479, 
    6196, 
    4845, 
    6201, 
    4997, 
    5140, 
    5941, 
    5609, 
    5337, 
    3337, 
    6114, 
    5609, 
    4086, 
    1142, 
    6114, 
    4086, 
    1378, 
    1622, 
    6114, 
    2590, 
    5337, 
    5609, 
    4086, 
    3001, 
    1142, 
    5912, 
    4995, 
    1461, 
    1879, 
    5912, 
    1052, 
    5704, 
    4995, 
    5912, 
    2642, 
    5704, 
    3001, 
    2642, 
    6002, 
    5704, 
    5704, 
    5912, 
    1879, 
    2400, 
    5021, 
    1714, 
    1879, 
    1345, 
    1142, 
    4579, 
    5965, 
    4386, 
    6114, 
    2329, 
    1378, 
    2400, 
    870, 
    1251, 
    6503, 
    4699, 
    6195, 
    5253, 
    5140, 
    5918, 
    3807, 
    5253, 
    5021, 
    3807, 
    3528, 
    5847, 
    5847, 
    3528, 
    5807, 
    5941, 
    5847, 
    5807, 
    5253, 
    3807, 
    5847, 
    1251, 
    3807, 
    2400, 
    5445, 
    5918, 
    4997, 
    5613, 
    2329, 
    4527, 
    4699, 
    5613, 
    4527, 
    5445, 
    1019, 
    6149, 
    6015, 
    921, 
    1714, 
    6503, 
    3931, 
    3658, 
    4871, 
    6503, 
    5023, 
    6195, 
    3931, 
    6503, 
    1345, 
    4171, 
    4527, 
    1345, 
    1052, 
    5965, 
    4579, 
    3931, 
    4171, 
    4584, 
    4579, 
    4386, 
    1548, 
    700, 
    5293, 
    1633, 
    1424, 
    5475, 
    3658, 
    3931, 
    4579, 
    5188, 
    2803, 
    4913, 
    3070, 
    6327, 
    4913, 
    921, 
    2068, 
    5188, 
    6008, 
    1756, 
    5871, 
    2922, 
    6008, 
    2511, 
    1560, 
    1756, 
    6008, 
    277, 
    1210, 
    278, 
    276, 
    275, 
    1800, 
    1798, 
    5736, 
    2358, 
    5114, 
    1558, 
    4250, 
    4460, 
    5114, 
    4250, 
    2984, 
    2593, 
    5114, 
    1033, 
    2984, 
    1798, 
    2593, 
    717, 
    5114, 
    845, 
    731, 
    1731, 
    6251, 
    1216, 
    947, 
    2370, 
    3471, 
    1418, 
    5840, 
    6363, 
    2899, 
    6251, 
    5888, 
    2792, 
    2370, 
    1849, 
    6363, 
    1558, 
    2370, 
    1418, 
    3471, 
    5840, 
    2792, 
    4978, 
    5871, 
    1756, 
    2291, 
    4978, 
    1756, 
    1800, 
    847, 
    5218, 
    3143, 
    4802, 
    4956, 
    870, 
    3070, 
    4629, 
    870, 
    1714, 
    6327, 
    4802, 
    4629, 
    3070, 
    5438, 
    4956, 
    2694, 
    3143, 
    3465, 
    4802, 
    1731, 
    2277, 
    5281, 
    5438, 
    1274, 
    4197, 
    5438, 
    1973, 
    1274, 
    4913, 
    3965, 
    2694, 
    3158, 
    746, 
    3965, 
    746, 
    3478, 
    3744, 
    3744, 
    1835, 
    1081, 
    1973, 
    3744, 
    1274, 
    1973, 
    746, 
    3744, 
    5823, 
    881, 
    1687, 
    5710, 
    1187, 
    2387, 
    3925, 
    5962, 
    2387, 
    4905, 
    2662, 
    5710, 
    731, 
    1964, 
    945, 
    4795, 
    1392, 
    1964, 
    731, 
    4795, 
    1964, 
    731, 
    4111, 
    4795, 
    4111, 
    731, 
    845, 
    3844, 
    4111, 
    845, 
    2353, 
    4795, 
    4111, 
    1330, 
    706, 
    1550, 
    4920, 
    1330, 
    1105, 
    4295, 
    1238, 
    2850, 
    1288, 
    758, 
    904, 
    1486, 
    1288, 
    904, 
    1002, 
    1486, 
    904, 
    1002, 
    756, 
    2850, 
    1238, 
    1743, 
    2285, 
    2253, 
    1238, 
    2285, 
    1486, 
    2253, 
    1288, 
    1486, 
    1002, 
    2850, 
    1171, 
    957, 
    1743, 
    1704, 
    3928, 
    209, 
    2850, 
    1238, 
    2253, 
    1486, 
    2850, 
    2253, 
    756, 
    1591, 
    2850, 
    758, 
    211, 
    904, 
    3694, 
    1221, 
    2240, 
    6240, 
    3097, 
    3694, 
    6250, 
    6240, 
    3400, 
    3425, 
    3097, 
    6240, 
    2689, 
    6143, 
    6250, 
    2507, 
    2919, 
    4424, 
    4424, 
    2919, 
    677, 
    3425, 
    4424, 
    3097, 
    3425, 
    2507, 
    4424, 
    1696, 
    2247, 
    677, 
    1233, 
    1221, 
    1936, 
    4612, 
    2142, 
    2571, 
    1844, 
    4612, 
    2571, 
    3048, 
    2666, 
    4612, 
    1943, 
    1221, 
    1233, 
    1046, 
    205, 
    2136, 
    4280, 
    5993, 
    6218, 
    2136, 
    4059, 
    1046, 
    2136, 
    1544, 
    4059, 
    206, 
    205, 
    1046, 
    4231, 
    6153, 
    2046, 
    5183, 
    6223, 
    1612, 
    6536, 
    6085, 
    6202, 
    5973, 
    6536, 
    5760, 
    5973, 
    6085, 
    6536, 
    4905, 
    5710, 
    5962, 
    5760, 
    4905, 
    5049, 
    2662, 
    1964, 
    5710, 
    881, 
    2387, 
    1187, 
    5183, 
    1612, 
    778, 
    1129, 
    3653, 
    3925, 
    1129, 
    288, 
    3653, 
    1956, 
    1100, 
    1849, 
    2593, 
    1956, 
    717, 
    1558, 
    5114, 
    717, 
    5757, 
    1033, 
    5322, 
    5225, 
    5757, 
    5322, 
    2984, 
    1033, 
    5757, 
    1250, 
    1100, 
    1956, 
    5322, 
    4330, 
    4530, 
    4330, 
    1535, 
    2919, 
    1250, 
    1956, 
    5225, 
    2129, 
    1535, 
    4330, 
    2052, 
    2129, 
    1033, 
    2052, 
    895, 
    2129, 
    6406, 
    2507, 
    3717, 
    919, 
    6406, 
    3717, 
    6246, 
    2507, 
    6406, 
    4530, 
    6246, 
    2263, 
    4530, 
    5731, 
    6246, 
    1250, 
    4530, 
    2263, 
    4330, 
    5731, 
    4530, 
    2263, 
    2171, 
    1250, 
    2263, 
    1586, 
    2171, 
    5225, 
    5322, 
    4530, 
    1250, 
    5225, 
    4530, 
    2593, 
    2984, 
    5757, 
    6246, 
    6405, 
    2263, 
    6073, 
    3454, 
    3130, 
    3984, 
    5246, 
    4896, 
    5516, 
    3742, 
    3454, 
    752, 
    5516, 
    5246, 
    752, 
    919, 
    6226, 
    3996, 
    4066, 
    1552, 
    5018, 
    4732, 
    1951, 
    4732, 
    947, 
    4285, 
    5888, 
    1418, 
    3471, 
    2792, 
    5888, 
    3471, 
    5079, 
    1418, 
    5888, 
    877, 
    3727, 
    1683, 
    916, 
    1066, 
    2065, 
    1216, 
    1451, 
    4256, 
    1046, 
    207, 
    206, 
    1807, 
    207, 
    1046, 
    1046, 
    4059, 
    4280, 
    1393, 
    202, 
    612, 
    4808, 
    6290, 
    3592, 
    1824, 
    4631, 
    200, 
    1824, 
    4241, 
    5858, 
    4808, 
    3592, 
    2046, 
    4631, 
    4808, 
    1393, 
    4631, 
    5858, 
    6290, 
    6695, 
    204, 
    203, 
    202, 
    1113, 
    6695, 
    6695, 
    613, 
    204, 
    202, 
    6695, 
    203, 
    1113, 
    613, 
    6695, 
    2046, 
    1113, 
    202, 
    5368, 
    2046, 
    202, 
    1393, 
    5368, 
    202, 
    1393, 
    4808, 
    5368, 
    4231, 
    1544, 
    2136, 
    6153, 
    4231, 
    2136, 
    205, 
    6153, 
    2136, 
    1113, 
    2046, 
    6153, 
    884, 
    1544, 
    4231, 
    205, 
    613, 
    1113, 
    1107, 
    1824, 
    199, 
    1453, 
    1069, 
    192, 
    1453, 
    1104, 
    4012, 
    5762, 
    4406, 
    1453, 
    191, 
    5762, 
    192, 
    191, 
    1741, 
    5762, 
    5799, 
    3961, 
    4192, 
    4408, 
    5986, 
    6179, 
    4605, 
    4406, 
    5799, 
    192, 
    5762, 
    1453, 
    997, 
    3961, 
    4406, 
    5858, 
    4241, 
    4012, 
    949, 
    2541, 
    1104, 
    949, 
    1737, 
    4607, 
    1824, 
    200, 
    199, 
    1453, 
    4012, 
    1069, 
    5100, 
    2541, 
    2946, 
    5858, 
    5100, 
    2946, 
    3286, 
    6290, 
    2946, 
    4631, 
    1824, 
    5858, 
    4012, 
    1104, 
    5100, 
    3097, 
    1936, 
    1221, 
    6405, 
    6246, 
    6406, 
    752, 
    6405, 
    919, 
    752, 
    1586, 
    6405, 
    4424, 
    1936, 
    3097, 
    5731, 
    2919, 
    2507, 
    6246, 
    5731, 
    2507, 
    4330, 
    2919, 
    5731, 
    677, 
    1936, 
    4424, 
    6153, 
    205, 
    1113, 
    884, 
    4231, 
    2046, 
    1544, 
    2775, 
    5993, 
    1689, 
    1544, 
    884, 
    692, 
    2600, 
    2775, 
    1393, 
    201, 
    200, 
    1393, 
    612, 
    201, 
    1350, 
    197, 
    196, 
    1350, 
    611, 
    198, 
    197, 
    1350, 
    198, 
    196, 
    610, 
    3207, 
    3207, 
    610, 
    6595, 
    6595, 
    610, 
    195, 
    194, 
    6595, 
    195, 
    194, 
    3207, 
    6595, 
    3207, 
    1286, 
    611, 
    196, 
    3207, 
    1350, 
    194, 
    1286, 
    3207, 
    3207, 
    611, 
    1350, 
    193, 
    1286, 
    194, 
    199, 
    611, 
    1286, 
    1107, 
    1286, 
    193, 
    1069, 
    193, 
    192, 
    1107, 
    199, 
    1286, 
    1069, 
    1107, 
    193, 
    1069, 
    1824, 
    1107, 
    3720, 
    670, 
    1529, 
    2144, 
    3429, 
    1060, 
    1451, 
    670, 
    3429, 
    2144, 
    4256, 
    3429, 
    5305, 
    3220, 
    2750, 
    1817, 
    2870, 
    1060, 
    1817, 
    2913, 
    4982, 
    1552, 
    4256, 
    2144, 
    1216, 
    6088, 
    1451, 
    5079, 
    2065, 
    1418, 
    6251, 
    5079, 
    5888, 
    1216, 
    6251, 
    2792, 
    1683, 
    5079, 
    6251, 
    1683, 
    3727, 
    5079, 
    1734, 
    1683, 
    947, 
    4285, 
    709, 
    4732, 
    5833, 
    4285, 
    947, 
    1216, 
    5833, 
    947, 
    4256, 
    1552, 
    5833, 
    709, 
    1951, 
    4732, 
    5018, 
    3681, 
    1277, 
    4732, 
    5018, 
    2280, 
    1244, 
    3681, 
    5018, 
    5079, 
    3727, 
    2065, 
    2792, 
    5840, 
    6088, 
    2593, 
    5225, 
    1956, 
    2483, 
    3099, 
    670, 
    1250, 
    2171, 
    1100, 
    3099, 
    1529, 
    670, 
    3427, 
    3099, 
    2483, 
    3718, 
    3427, 
    2899, 
    1100, 
    3718, 
    2899, 
    2171, 
    1586, 
    3984, 
    3718, 
    2171, 
    3984, 
    5246, 
    3984, 
    1586, 
    1027, 
    6310, 
    2767, 
    6315, 
    3984, 
    4896, 
    4607, 
    1422, 
    2689, 
    1535, 
    1696, 
    677, 
    692, 
    1544, 
    1689, 
    5645, 
    3706, 
    4192, 
    5100, 
    1104, 
    2541, 
    6290, 
    4808, 
    4631, 
    2946, 
    6290, 
    5858, 
    3286, 
    3592, 
    6290, 
    4241, 
    1069, 
    4012, 
    5100, 
    5858, 
    4012, 
    1824, 
    1069, 
    4241, 
    3717, 
    6143, 
    919, 
    3694, 
    3395, 
    4193, 
    6240, 
    3694, 
    3400, 
    2240, 
    3395, 
    3694, 
    3694, 
    3097, 
    1221, 
    4193, 
    3400, 
    3694, 
    3286, 
    4193, 
    3395, 
    3286, 
    2946, 
    4193, 
    6143, 
    1422, 
    1280, 
    3425, 
    6250, 
    3717, 
    2689, 
    1422, 
    6143, 
    1943, 
    2240, 
    1221, 
    1943, 
    692, 
    2240, 
    4607, 
    2541, 
    949, 
    1422, 
    4607, 
    1737, 
    4409, 
    2541, 
    4607, 
    3400, 
    4193, 
    4409, 
    3592, 
    3286, 
    3395, 
    1689, 
    3592, 
    3395, 
    884, 
    2046, 
    3592, 
    4808, 
    2046, 
    5368, 
    4631, 
    1393, 
    200, 
    2689, 
    4409, 
    4607, 
    1280, 
    919, 
    6143, 
    3592, 
    1689, 
    884, 
    4409, 
    2689, 
    3400, 
    2946, 
    4409, 
    4193, 
    2946, 
    2541, 
    4409, 
    2240, 
    1689, 
    3395, 
    5762, 
    997, 
    4406, 
    4827, 
    3130, 
    4649, 
    6060, 
    4827, 
    4649, 
    4980, 
    781, 
    1615, 
    4683, 
    4980, 
    4827, 
    4683, 
    1357, 
    4980, 
    6405, 
    1586, 
    2263, 
    5450, 
    4827, 
    4980, 
    6250, 
    3425, 
    6240, 
    2689, 
    6250, 
    3400, 
    6143, 
    3717, 
    6250, 
    6405, 
    6406, 
    919, 
    2507, 
    3425, 
    3717, 
    1357, 
    4683, 
    6392, 
    6121, 
    4649, 
    3742, 
    6524, 
    6121, 
    5626, 
    3693, 
    6524, 
    5626, 
    4298, 
    6121, 
    6524, 
    4298, 
    6060, 
    6121, 
    6073, 
    5516, 
    3454, 
    6226, 
    1280, 
    3742, 
    184, 
    609, 
    2704, 
    1626, 
    797, 
    1088, 
    1145, 
    5503, 
    1037, 
    5066, 
    3238, 
    3549, 
    5005, 
    666, 
    982, 
    3409, 
    5005, 
    982, 
    3706, 
    2704, 
    5005 ;

 grid.cells.vertex_refs_start = 
    0, 
    3, 
    6, 
    9, 
    12, 
    15, 
    18, 
    21, 
    24, 
    27, 
    30, 
    33, 
    36, 
    39, 
    42, 
    45, 
    48, 
    51, 
    54, 
    57, 
    60, 
    63, 
    66, 
    69, 
    72, 
    75, 
    78, 
    81, 
    84, 
    87, 
    90, 
    93, 
    96, 
    99, 
    102, 
    105, 
    108, 
    111, 
    114, 
    117, 
    120, 
    123, 
    126, 
    129, 
    132, 
    135, 
    138, 
    141, 
    144, 
    147, 
    150, 
    153, 
    156, 
    159, 
    162, 
    165, 
    168, 
    171, 
    174, 
    177, 
    180, 
    183, 
    186, 
    189, 
    192, 
    195, 
    198, 
    201, 
    204, 
    207, 
    210, 
    213, 
    216, 
    219, 
    222, 
    225, 
    228, 
    231, 
    234, 
    237, 
    240, 
    243, 
    246, 
    249, 
    252, 
    255, 
    258, 
    261, 
    264, 
    267, 
    270, 
    273, 
    276, 
    279, 
    282, 
    285, 
    288, 
    291, 
    294, 
    297, 
    300, 
    303, 
    306, 
    309, 
    312, 
    315, 
    318, 
    321, 
    324, 
    327, 
    330, 
    333, 
    336, 
    339, 
    342, 
    345, 
    348, 
    351, 
    354, 
    357, 
    360, 
    363, 
    366, 
    369, 
    372, 
    375, 
    378, 
    381, 
    384, 
    387, 
    390, 
    393, 
    396, 
    399, 
    402, 
    405, 
    408, 
    411, 
    414, 
    417, 
    420, 
    423, 
    426, 
    429, 
    432, 
    435, 
    438, 
    441, 
    444, 
    447, 
    450, 
    453, 
    456, 
    459, 
    462, 
    465, 
    468, 
    471, 
    474, 
    477, 
    480, 
    483, 
    486, 
    489, 
    492, 
    495, 
    498, 
    501, 
    504, 
    507, 
    510, 
    513, 
    516, 
    519, 
    522, 
    525, 
    528, 
    531, 
    534, 
    537, 
    540, 
    543, 
    546, 
    549, 
    552, 
    555, 
    558, 
    561, 
    564, 
    567, 
    570, 
    573, 
    576, 
    579, 
    582, 
    585, 
    588, 
    591, 
    594, 
    597, 
    600, 
    603, 
    606, 
    609, 
    612, 
    615, 
    618, 
    621, 
    624, 
    627, 
    630, 
    633, 
    636, 
    639, 
    642, 
    645, 
    648, 
    651, 
    654, 
    657, 
    660, 
    663, 
    666, 
    669, 
    672, 
    675, 
    678, 
    681, 
    684, 
    687, 
    690, 
    693, 
    696, 
    699, 
    702, 
    705, 
    708, 
    711, 
    714, 
    717, 
    720, 
    723, 
    726, 
    729, 
    732, 
    735, 
    738, 
    741, 
    744, 
    747, 
    750, 
    753, 
    756, 
    759, 
    762, 
    765, 
    768, 
    771, 
    774, 
    777, 
    780, 
    783, 
    786, 
    789, 
    792, 
    795, 
    798, 
    801, 
    804, 
    807, 
    810, 
    813, 
    816, 
    819, 
    822, 
    825, 
    828, 
    831, 
    834, 
    837, 
    840, 
    843, 
    846, 
    849, 
    852, 
    855, 
    858, 
    861, 
    864, 
    867, 
    870, 
    873, 
    876, 
    879, 
    882, 
    885, 
    888, 
    891, 
    894, 
    897, 
    900, 
    903, 
    906, 
    909, 
    912, 
    915, 
    918, 
    921, 
    924, 
    927, 
    930, 
    933, 
    936, 
    939, 
    942, 
    945, 
    948, 
    951, 
    954, 
    957, 
    960, 
    963, 
    966, 
    969, 
    972, 
    975, 
    978, 
    981, 
    984, 
    987, 
    990, 
    993, 
    996, 
    999, 
    1002, 
    1005, 
    1008, 
    1011, 
    1014, 
    1017, 
    1020, 
    1023, 
    1026, 
    1029, 
    1032, 
    1035, 
    1038, 
    1041, 
    1044, 
    1047, 
    1050, 
    1053, 
    1056, 
    1059, 
    1062, 
    1065, 
    1068, 
    1071, 
    1074, 
    1077, 
    1080, 
    1083, 
    1086, 
    1089, 
    1092, 
    1095, 
    1098, 
    1101, 
    1104, 
    1107, 
    1110, 
    1113, 
    1116, 
    1119, 
    1122, 
    1125, 
    1128, 
    1131, 
    1134, 
    1137, 
    1140, 
    1143, 
    1146, 
    1149, 
    1152, 
    1155, 
    1158, 
    1161, 
    1164, 
    1167, 
    1170, 
    1173, 
    1176, 
    1179, 
    1182, 
    1185, 
    1188, 
    1191, 
    1194, 
    1197, 
    1200, 
    1203, 
    1206, 
    1209, 
    1212, 
    1215, 
    1218, 
    1221, 
    1224, 
    1227, 
    1230, 
    1233, 
    1236, 
    1239, 
    1242, 
    1245, 
    1248, 
    1251, 
    1254, 
    1257, 
    1260, 
    1263, 
    1266, 
    1269, 
    1272, 
    1275, 
    1278, 
    1281, 
    1284, 
    1287, 
    1290, 
    1293, 
    1296, 
    1299, 
    1302, 
    1305, 
    1308, 
    1311, 
    1314, 
    1317, 
    1320, 
    1323, 
    1326, 
    1329, 
    1332, 
    1335, 
    1338, 
    1341, 
    1344, 
    1347, 
    1350, 
    1353, 
    1356, 
    1359, 
    1362, 
    1365, 
    1368, 
    1371, 
    1374, 
    1377, 
    1380, 
    1383, 
    1386, 
    1389, 
    1392, 
    1395, 
    1398, 
    1401, 
    1404, 
    1407, 
    1410, 
    1413, 
    1416, 
    1419, 
    1422, 
    1425, 
    1428, 
    1431, 
    1434, 
    1437, 
    1440, 
    1443, 
    1446, 
    1449, 
    1452, 
    1455, 
    1458, 
    1461, 
    1464, 
    1467, 
    1470, 
    1473, 
    1476, 
    1479, 
    1482, 
    1485, 
    1488, 
    1491, 
    1494, 
    1497, 
    1500, 
    1503, 
    1506, 
    1509, 
    1512, 
    1515, 
    1518, 
    1521, 
    1524, 
    1527, 
    1530, 
    1533, 
    1536, 
    1539, 
    1542, 
    1545, 
    1548, 
    1551, 
    1554, 
    1557, 
    1560, 
    1563, 
    1566, 
    1569, 
    1572, 
    1575, 
    1578, 
    1581, 
    1584, 
    1587, 
    1590, 
    1593, 
    1596, 
    1599, 
    1602, 
    1605, 
    1608, 
    1611, 
    1614, 
    1617, 
    1620, 
    1623, 
    1626, 
    1629, 
    1632, 
    1635, 
    1638, 
    1641, 
    1644, 
    1647, 
    1650, 
    1653, 
    1656, 
    1659, 
    1662, 
    1665, 
    1668, 
    1671, 
    1674, 
    1677, 
    1680, 
    1683, 
    1686, 
    1689, 
    1692, 
    1695, 
    1698, 
    1701, 
    1704, 
    1707, 
    1710, 
    1713, 
    1716, 
    1719, 
    1722, 
    1725, 
    1728, 
    1731, 
    1734, 
    1737, 
    1740, 
    1743, 
    1746, 
    1749, 
    1752, 
    1755, 
    1758, 
    1761, 
    1764, 
    1767, 
    1770, 
    1773, 
    1776, 
    1779, 
    1782, 
    1785, 
    1788, 
    1791, 
    1794, 
    1797, 
    1800, 
    1803, 
    1806, 
    1809, 
    1812, 
    1815, 
    1818, 
    1821, 
    1824, 
    1827, 
    1830, 
    1833, 
    1836, 
    1839, 
    1842, 
    1845, 
    1848, 
    1851, 
    1854, 
    1857, 
    1860, 
    1863, 
    1866, 
    1869, 
    1872, 
    1875, 
    1878, 
    1881, 
    1884, 
    1887, 
    1890, 
    1893, 
    1896, 
    1899, 
    1902, 
    1905, 
    1908, 
    1911, 
    1914, 
    1917, 
    1920, 
    1923, 
    1926, 
    1929, 
    1932, 
    1935, 
    1938, 
    1941, 
    1944, 
    1947, 
    1950, 
    1953, 
    1956, 
    1959, 
    1962, 
    1965, 
    1968, 
    1971, 
    1974, 
    1977, 
    1980, 
    1983, 
    1986, 
    1989, 
    1992, 
    1995, 
    1998, 
    2001, 
    2004, 
    2007, 
    2010, 
    2013, 
    2016, 
    2019, 
    2022, 
    2025, 
    2028, 
    2031, 
    2034, 
    2037, 
    2040, 
    2043, 
    2046, 
    2049, 
    2052, 
    2055, 
    2058, 
    2061, 
    2064, 
    2067, 
    2070, 
    2073, 
    2076, 
    2079, 
    2082, 
    2085, 
    2088, 
    2091, 
    2094, 
    2097, 
    2100, 
    2103, 
    2106, 
    2109, 
    2112, 
    2115, 
    2118, 
    2121, 
    2124, 
    2127, 
    2130, 
    2133, 
    2136, 
    2139, 
    2142, 
    2145, 
    2148, 
    2151, 
    2154, 
    2157, 
    2160, 
    2163, 
    2166, 
    2169, 
    2172, 
    2175, 
    2178, 
    2181, 
    2184, 
    2187, 
    2190, 
    2193, 
    2196, 
    2199, 
    2202, 
    2205, 
    2208, 
    2211, 
    2214, 
    2217, 
    2220, 
    2223, 
    2226, 
    2229, 
    2232, 
    2235, 
    2238, 
    2241, 
    2244, 
    2247, 
    2250, 
    2253, 
    2256, 
    2259, 
    2262, 
    2265, 
    2268, 
    2271, 
    2274, 
    2277, 
    2280, 
    2283, 
    2286, 
    2289, 
    2292, 
    2295, 
    2298, 
    2301, 
    2304, 
    2307, 
    2310, 
    2313, 
    2316, 
    2319, 
    2322, 
    2325, 
    2328, 
    2331, 
    2334, 
    2337, 
    2340, 
    2343, 
    2346, 
    2349, 
    2352, 
    2355, 
    2358, 
    2361, 
    2364, 
    2367, 
    2370, 
    2373, 
    2376, 
    2379, 
    2382, 
    2385, 
    2388, 
    2391, 
    2394, 
    2397, 
    2400, 
    2403, 
    2406, 
    2409, 
    2412, 
    2415, 
    2418, 
    2421, 
    2424, 
    2427, 
    2430, 
    2433, 
    2436, 
    2439, 
    2442, 
    2445, 
    2448, 
    2451, 
    2454, 
    2457, 
    2460, 
    2463, 
    2466, 
    2469, 
    2472, 
    2475, 
    2478, 
    2481, 
    2484, 
    2487, 
    2490, 
    2493, 
    2496, 
    2499, 
    2502, 
    2505, 
    2508, 
    2511, 
    2514, 
    2517, 
    2520, 
    2523, 
    2526, 
    2529, 
    2532, 
    2535, 
    2538, 
    2541, 
    2544, 
    2547, 
    2550, 
    2553, 
    2556, 
    2559, 
    2562, 
    2565, 
    2568, 
    2571, 
    2574, 
    2577, 
    2580, 
    2583, 
    2586, 
    2589, 
    2592, 
    2595, 
    2598, 
    2601, 
    2604, 
    2607, 
    2610, 
    2613, 
    2616, 
    2619, 
    2622, 
    2625, 
    2628, 
    2631, 
    2634, 
    2637, 
    2640, 
    2643, 
    2646, 
    2649, 
    2652, 
    2655, 
    2658, 
    2661, 
    2664, 
    2667, 
    2670, 
    2673, 
    2676, 
    2679, 
    2682, 
    2685, 
    2688, 
    2691, 
    2694, 
    2697, 
    2700, 
    2703, 
    2706, 
    2709, 
    2712, 
    2715, 
    2718, 
    2721, 
    2724, 
    2727, 
    2730, 
    2733, 
    2736, 
    2739, 
    2742, 
    2745, 
    2748, 
    2751, 
    2754, 
    2757, 
    2760, 
    2763, 
    2766, 
    2769, 
    2772, 
    2775, 
    2778, 
    2781, 
    2784, 
    2787, 
    2790, 
    2793, 
    2796, 
    2799, 
    2802, 
    2805, 
    2808, 
    2811, 
    2814, 
    2817, 
    2820, 
    2823, 
    2826, 
    2829, 
    2832, 
    2835, 
    2838, 
    2841, 
    2844, 
    2847, 
    2850, 
    2853, 
    2856, 
    2859, 
    2862, 
    2865, 
    2868, 
    2871, 
    2874, 
    2877, 
    2880, 
    2883, 
    2886, 
    2889, 
    2892, 
    2895, 
    2898, 
    2901, 
    2904, 
    2907, 
    2910, 
    2913, 
    2916, 
    2919, 
    2922, 
    2925, 
    2928, 
    2931, 
    2934, 
    2937, 
    2940, 
    2943, 
    2946, 
    2949, 
    2952, 
    2955, 
    2958, 
    2961, 
    2964, 
    2967, 
    2970, 
    2973, 
    2976, 
    2979, 
    2982, 
    2985, 
    2988, 
    2991, 
    2994, 
    2997, 
    3000, 
    3003, 
    3006, 
    3009, 
    3012, 
    3015, 
    3018, 
    3021, 
    3024, 
    3027, 
    3030, 
    3033, 
    3036, 
    3039, 
    3042, 
    3045, 
    3048, 
    3051, 
    3054, 
    3057, 
    3060, 
    3063, 
    3066, 
    3069, 
    3072, 
    3075, 
    3078, 
    3081, 
    3084, 
    3087, 
    3090, 
    3093, 
    3096, 
    3099, 
    3102, 
    3105, 
    3108, 
    3111, 
    3114, 
    3117, 
    3120, 
    3123, 
    3126, 
    3129, 
    3132, 
    3135, 
    3138, 
    3141, 
    3144, 
    3147, 
    3150, 
    3153, 
    3156, 
    3159, 
    3162, 
    3165, 
    3168, 
    3171, 
    3174, 
    3177, 
    3180, 
    3183, 
    3186, 
    3189, 
    3192, 
    3195, 
    3198, 
    3201, 
    3204, 
    3207, 
    3210, 
    3213, 
    3216, 
    3219, 
    3222, 
    3225, 
    3228, 
    3231, 
    3234, 
    3237, 
    3240, 
    3243, 
    3246, 
    3249, 
    3252, 
    3255, 
    3258, 
    3261, 
    3264, 
    3267, 
    3270, 
    3273, 
    3276, 
    3279, 
    3282, 
    3285, 
    3288, 
    3291, 
    3294, 
    3297, 
    3300, 
    3303, 
    3306, 
    3309, 
    3312, 
    3315, 
    3318, 
    3321, 
    3324, 
    3327, 
    3330, 
    3333, 
    3336, 
    3339, 
    3342, 
    3345, 
    3348, 
    3351, 
    3354, 
    3357, 
    3360, 
    3363, 
    3366, 
    3369, 
    3372, 
    3375, 
    3378, 
    3381, 
    3384, 
    3387, 
    3390, 
    3393, 
    3396, 
    3399, 
    3402, 
    3405, 
    3408, 
    3411, 
    3414, 
    3417, 
    3420, 
    3423, 
    3426, 
    3429, 
    3432, 
    3435, 
    3438, 
    3441, 
    3444, 
    3447, 
    3450, 
    3453, 
    3456, 
    3459, 
    3462, 
    3465, 
    3468, 
    3471, 
    3474, 
    3477, 
    3480, 
    3483, 
    3486, 
    3489, 
    3492, 
    3495, 
    3498, 
    3501, 
    3504, 
    3507, 
    3510, 
    3513, 
    3516, 
    3519, 
    3522, 
    3525, 
    3528, 
    3531, 
    3534, 
    3537, 
    3540, 
    3543, 
    3546, 
    3549, 
    3552, 
    3555, 
    3558, 
    3561, 
    3564, 
    3567, 
    3570, 
    3573, 
    3576, 
    3579, 
    3582, 
    3585, 
    3588, 
    3591, 
    3594, 
    3597, 
    3600, 
    3603, 
    3606, 
    3609, 
    3612, 
    3615, 
    3618, 
    3621, 
    3624, 
    3627, 
    3630, 
    3633, 
    3636, 
    3639, 
    3642, 
    3645, 
    3648, 
    3651, 
    3654, 
    3657, 
    3660, 
    3663, 
    3666, 
    3669, 
    3672, 
    3675, 
    3678, 
    3681, 
    3684, 
    3687, 
    3690, 
    3693, 
    3696, 
    3699, 
    3702, 
    3705, 
    3708, 
    3711, 
    3714, 
    3717, 
    3720, 
    3723, 
    3726, 
    3729, 
    3732, 
    3735, 
    3738, 
    3741, 
    3744, 
    3747, 
    3750, 
    3753, 
    3756, 
    3759, 
    3762, 
    3765, 
    3768, 
    3771, 
    3774, 
    3777, 
    3780, 
    3783, 
    3786, 
    3789, 
    3792, 
    3795, 
    3798, 
    3801, 
    3804, 
    3807, 
    3810, 
    3813, 
    3816, 
    3819, 
    3822, 
    3825, 
    3828, 
    3831, 
    3834, 
    3837, 
    3840, 
    3843, 
    3846, 
    3849, 
    3852, 
    3855, 
    3858, 
    3861, 
    3864, 
    3867, 
    3870, 
    3873, 
    3876, 
    3879, 
    3882, 
    3885, 
    3888, 
    3891, 
    3894, 
    3897, 
    3900, 
    3903, 
    3906, 
    3909, 
    3912, 
    3915, 
    3918, 
    3921, 
    3924, 
    3927, 
    3930, 
    3933, 
    3936, 
    3939, 
    3942, 
    3945, 
    3948, 
    3951, 
    3954, 
    3957, 
    3960, 
    3963, 
    3966, 
    3969, 
    3972, 
    3975, 
    3978, 
    3981, 
    3984, 
    3987, 
    3990, 
    3993, 
    3996, 
    3999, 
    4002, 
    4005, 
    4008, 
    4011, 
    4014, 
    4017, 
    4020, 
    4023, 
    4026, 
    4029, 
    4032, 
    4035, 
    4038, 
    4041, 
    4044, 
    4047, 
    4050, 
    4053, 
    4056, 
    4059, 
    4062, 
    4065, 
    4068, 
    4071, 
    4074, 
    4077, 
    4080, 
    4083, 
    4086, 
    4089, 
    4092, 
    4095, 
    4098, 
    4101, 
    4104, 
    4107, 
    4110, 
    4113, 
    4116, 
    4119, 
    4122, 
    4125, 
    4128, 
    4131, 
    4134, 
    4137, 
    4140, 
    4143, 
    4146, 
    4149, 
    4152, 
    4155, 
    4158, 
    4161, 
    4164, 
    4167, 
    4170, 
    4173, 
    4176, 
    4179, 
    4182, 
    4185, 
    4188, 
    4191, 
    4194, 
    4197, 
    4200, 
    4203, 
    4206, 
    4209, 
    4212, 
    4215, 
    4218, 
    4221, 
    4224, 
    4227, 
    4230, 
    4233, 
    4236, 
    4239, 
    4242, 
    4245, 
    4248, 
    4251, 
    4254, 
    4257, 
    4260, 
    4263, 
    4266, 
    4269, 
    4272, 
    4275, 
    4278, 
    4281, 
    4284, 
    4287, 
    4290, 
    4293, 
    4296, 
    4299, 
    4302, 
    4305, 
    4308, 
    4311, 
    4314, 
    4317, 
    4320, 
    4323, 
    4326, 
    4329, 
    4332, 
    4335, 
    4338, 
    4341, 
    4344, 
    4347, 
    4350, 
    4353, 
    4356, 
    4359, 
    4362, 
    4365, 
    4368, 
    4371, 
    4374, 
    4377, 
    4380, 
    4383, 
    4386, 
    4389, 
    4392, 
    4395, 
    4398, 
    4401, 
    4404, 
    4407, 
    4410, 
    4413, 
    4416, 
    4419, 
    4422, 
    4425, 
    4428, 
    4431, 
    4434, 
    4437, 
    4440, 
    4443, 
    4446, 
    4449, 
    4452, 
    4455, 
    4458, 
    4461, 
    4464, 
    4467, 
    4470, 
    4473, 
    4476, 
    4479, 
    4482, 
    4485, 
    4488, 
    4491, 
    4494, 
    4497, 
    4500, 
    4503, 
    4506, 
    4509, 
    4512, 
    4515, 
    4518, 
    4521, 
    4524, 
    4527, 
    4530, 
    4533, 
    4536, 
    4539, 
    4542, 
    4545, 
    4548, 
    4551, 
    4554, 
    4557, 
    4560, 
    4563, 
    4566, 
    4569, 
    4572, 
    4575, 
    4578, 
    4581, 
    4584, 
    4587, 
    4590, 
    4593, 
    4596, 
    4599, 
    4602, 
    4605, 
    4608, 
    4611, 
    4614, 
    4617, 
    4620, 
    4623, 
    4626, 
    4629, 
    4632, 
    4635, 
    4638, 
    4641, 
    4644, 
    4647, 
    4650, 
    4653, 
    4656, 
    4659, 
    4662, 
    4665, 
    4668, 
    4671, 
    4674, 
    4677, 
    4680, 
    4683, 
    4686, 
    4689, 
    4692, 
    4695, 
    4698, 
    4701, 
    4704, 
    4707, 
    4710, 
    4713, 
    4716, 
    4719, 
    4722, 
    4725, 
    4728, 
    4731, 
    4734, 
    4737, 
    4740, 
    4743, 
    4746, 
    4749, 
    4752, 
    4755, 
    4758, 
    4761, 
    4764, 
    4767, 
    4770, 
    4773, 
    4776, 
    4779, 
    4782, 
    4785, 
    4788, 
    4791, 
    4794, 
    4797, 
    4800, 
    4803, 
    4806, 
    4809, 
    4812, 
    4815, 
    4818, 
    4821, 
    4824, 
    4827, 
    4830, 
    4833, 
    4836, 
    4839, 
    4842, 
    4845, 
    4848, 
    4851, 
    4854, 
    4857, 
    4860, 
    4863, 
    4866, 
    4869, 
    4872, 
    4875, 
    4878, 
    4881, 
    4884, 
    4887, 
    4890, 
    4893, 
    4896, 
    4899, 
    4902, 
    4905, 
    4908, 
    4911, 
    4914, 
    4917, 
    4920, 
    4923, 
    4926, 
    4929, 
    4932, 
    4935, 
    4938, 
    4941, 
    4944, 
    4947, 
    4950, 
    4953, 
    4956, 
    4959, 
    4962, 
    4965, 
    4968, 
    4971, 
    4974, 
    4977, 
    4980, 
    4983, 
    4986, 
    4989, 
    4992, 
    4995, 
    4998, 
    5001, 
    5004, 
    5007, 
    5010, 
    5013, 
    5016, 
    5019, 
    5022, 
    5025, 
    5028, 
    5031, 
    5034, 
    5037, 
    5040, 
    5043, 
    5046, 
    5049, 
    5052, 
    5055, 
    5058, 
    5061, 
    5064, 
    5067, 
    5070, 
    5073, 
    5076, 
    5079, 
    5082, 
    5085, 
    5088, 
    5091, 
    5094, 
    5097, 
    5100, 
    5103, 
    5106, 
    5109, 
    5112, 
    5115, 
    5118, 
    5121, 
    5124, 
    5127, 
    5130, 
    5133, 
    5136, 
    5139, 
    5142, 
    5145, 
    5148, 
    5151, 
    5154, 
    5157, 
    5160, 
    5163, 
    5166, 
    5169, 
    5172, 
    5175, 
    5178, 
    5181, 
    5184, 
    5187, 
    5190, 
    5193, 
    5196, 
    5199, 
    5202, 
    5205, 
    5208, 
    5211, 
    5214, 
    5217, 
    5220, 
    5223, 
    5226, 
    5229, 
    5232, 
    5235, 
    5238, 
    5241, 
    5244, 
    5247, 
    5250, 
    5253, 
    5256, 
    5259, 
    5262, 
    5265, 
    5268, 
    5271, 
    5274, 
    5277, 
    5280, 
    5283, 
    5286, 
    5289, 
    5292, 
    5295, 
    5298, 
    5301, 
    5304, 
    5307, 
    5310, 
    5313, 
    5316, 
    5319, 
    5322, 
    5325, 
    5328, 
    5331, 
    5334, 
    5337, 
    5340, 
    5343, 
    5346, 
    5349, 
    5352, 
    5355, 
    5358, 
    5361, 
    5364, 
    5367, 
    5370, 
    5373, 
    5376, 
    5379, 
    5382, 
    5385, 
    5388, 
    5391, 
    5394, 
    5397, 
    5400, 
    5403, 
    5406, 
    5409, 
    5412, 
    5415, 
    5418, 
    5421, 
    5424, 
    5427, 
    5430, 
    5433, 
    5436, 
    5439, 
    5442, 
    5445, 
    5448, 
    5451, 
    5454, 
    5457, 
    5460, 
    5463, 
    5466, 
    5469, 
    5472, 
    5475, 
    5478, 
    5481, 
    5484, 
    5487, 
    5490, 
    5493, 
    5496, 
    5499, 
    5502, 
    5505, 
    5508, 
    5511, 
    5514, 
    5517, 
    5520, 
    5523, 
    5526, 
    5529, 
    5532, 
    5535, 
    5538, 
    5541, 
    5544, 
    5547, 
    5550, 
    5553, 
    5556, 
    5559, 
    5562, 
    5565, 
    5568, 
    5571, 
    5574, 
    5577, 
    5580, 
    5583, 
    5586, 
    5589, 
    5592, 
    5595, 
    5598, 
    5601, 
    5604, 
    5607, 
    5610, 
    5613, 
    5616, 
    5619, 
    5622, 
    5625, 
    5628, 
    5631, 
    5634, 
    5637, 
    5640, 
    5643, 
    5646, 
    5649, 
    5652, 
    5655, 
    5658, 
    5661, 
    5664, 
    5667, 
    5670, 
    5673, 
    5676, 
    5679, 
    5682, 
    5685, 
    5688, 
    5691, 
    5694, 
    5697, 
    5700, 
    5703, 
    5706, 
    5709, 
    5712, 
    5715, 
    5718, 
    5721, 
    5724, 
    5727, 
    5730, 
    5733, 
    5736, 
    5739, 
    5742, 
    5745, 
    5748, 
    5751, 
    5754, 
    5757, 
    5760, 
    5763, 
    5766, 
    5769, 
    5772, 
    5775, 
    5778, 
    5781, 
    5784, 
    5787, 
    5790, 
    5793, 
    5796, 
    5799, 
    5802, 
    5805, 
    5808, 
    5811, 
    5814, 
    5817, 
    5820, 
    5823, 
    5826, 
    5829, 
    5832, 
    5835, 
    5838, 
    5841, 
    5844, 
    5847, 
    5850, 
    5853, 
    5856, 
    5859, 
    5862, 
    5865, 
    5868, 
    5871, 
    5874, 
    5877, 
    5880, 
    5883, 
    5886, 
    5889, 
    5892, 
    5895, 
    5898, 
    5901, 
    5904, 
    5907, 
    5910, 
    5913, 
    5916, 
    5919, 
    5922, 
    5925, 
    5928, 
    5931, 
    5934, 
    5937, 
    5940, 
    5943, 
    5946, 
    5949, 
    5952, 
    5955, 
    5958, 
    5961, 
    5964, 
    5967, 
    5970, 
    5973, 
    5976, 
    5979, 
    5982, 
    5985, 
    5988, 
    5991, 
    5994, 
    5997, 
    6000, 
    6003, 
    6006, 
    6009, 
    6012, 
    6015, 
    6018, 
    6021, 
    6024, 
    6027, 
    6030, 
    6033, 
    6036, 
    6039, 
    6042, 
    6045, 
    6048, 
    6051, 
    6054, 
    6057, 
    6060, 
    6063, 
    6066, 
    6069, 
    6072, 
    6075, 
    6078, 
    6081, 
    6084, 
    6087, 
    6090, 
    6093, 
    6096, 
    6099, 
    6102, 
    6105, 
    6108, 
    6111, 
    6114, 
    6117, 
    6120, 
    6123, 
    6126, 
    6129, 
    6132, 
    6135, 
    6138, 
    6141, 
    6144, 
    6147, 
    6150, 
    6153, 
    6156, 
    6159, 
    6162, 
    6165, 
    6168, 
    6171, 
    6174, 
    6177, 
    6180, 
    6183, 
    6186, 
    6189, 
    6192, 
    6195, 
    6198, 
    6201, 
    6204, 
    6207, 
    6210, 
    6213, 
    6216, 
    6219, 
    6222, 
    6225, 
    6228, 
    6231, 
    6234, 
    6237, 
    6240, 
    6243, 
    6246, 
    6249, 
    6252, 
    6255, 
    6258, 
    6261, 
    6264, 
    6267, 
    6270, 
    6273, 
    6276, 
    6279, 
    6282, 
    6285, 
    6288, 
    6291, 
    6294, 
    6297, 
    6300, 
    6303, 
    6306, 
    6309, 
    6312, 
    6315, 
    6318, 
    6321, 
    6324, 
    6327, 
    6330, 
    6333, 
    6336, 
    6339, 
    6342, 
    6345, 
    6348, 
    6351, 
    6354, 
    6357, 
    6360, 
    6363, 
    6366, 
    6369, 
    6372, 
    6375, 
    6378, 
    6381, 
    6384, 
    6387, 
    6390, 
    6393, 
    6396, 
    6399, 
    6402, 
    6405, 
    6408, 
    6411, 
    6414, 
    6417, 
    6420, 
    6423, 
    6426, 
    6429, 
    6432, 
    6435, 
    6438, 
    6441, 
    6444, 
    6447, 
    6450, 
    6453, 
    6456, 
    6459, 
    6462, 
    6465, 
    6468, 
    6471, 
    6474, 
    6477, 
    6480, 
    6483, 
    6486, 
    6489, 
    6492, 
    6495, 
    6498, 
    6501, 
    6504, 
    6507, 
    6510, 
    6513, 
    6516, 
    6519, 
    6522, 
    6525, 
    6528, 
    6531, 
    6534, 
    6537, 
    6540, 
    6543, 
    6546, 
    6549, 
    6552, 
    6555, 
    6558, 
    6561, 
    6564, 
    6567, 
    6570, 
    6573, 
    6576, 
    6579, 
    6582, 
    6585, 
    6588, 
    6591, 
    6594, 
    6597, 
    6600, 
    6603, 
    6606, 
    6609, 
    6612, 
    6615, 
    6618, 
    6621, 
    6624, 
    6627, 
    6630, 
    6633, 
    6636, 
    6639, 
    6642, 
    6645, 
    6648, 
    6651, 
    6654, 
    6657, 
    6660, 
    6663, 
    6666, 
    6669, 
    6672, 
    6675, 
    6678, 
    6681, 
    6684, 
    6687, 
    6690, 
    6693, 
    6696, 
    6699, 
    6702, 
    6705, 
    6708, 
    6711, 
    6714, 
    6717, 
    6720, 
    6723, 
    6726, 
    6729, 
    6732, 
    6735, 
    6738, 
    6741, 
    6744, 
    6747, 
    6750, 
    6753, 
    6756, 
    6759, 
    6762, 
    6765, 
    6768, 
    6771, 
    6774, 
    6777, 
    6780, 
    6783, 
    6786, 
    6789, 
    6792, 
    6795, 
    6798, 
    6801, 
    6804, 
    6807, 
    6810, 
    6813, 
    6816, 
    6819, 
    6822, 
    6825, 
    6828, 
    6831, 
    6834, 
    6837, 
    6840, 
    6843, 
    6846, 
    6849, 
    6852, 
    6855, 
    6858, 
    6861, 
    6864, 
    6867, 
    6870, 
    6873, 
    6876, 
    6879, 
    6882, 
    6885, 
    6888, 
    6891, 
    6894, 
    6897, 
    6900, 
    6903, 
    6906, 
    6909, 
    6912, 
    6915, 
    6918, 
    6921, 
    6924, 
    6927, 
    6930, 
    6933, 
    6936, 
    6939, 
    6942, 
    6945, 
    6948, 
    6951, 
    6954, 
    6957, 
    6960, 
    6963, 
    6966, 
    6969, 
    6972, 
    6975, 
    6978, 
    6981, 
    6984, 
    6987, 
    6990, 
    6993, 
    6996, 
    6999, 
    7002, 
    7005, 
    7008, 
    7011, 
    7014, 
    7017, 
    7020, 
    7023, 
    7026, 
    7029, 
    7032, 
    7035, 
    7038, 
    7041, 
    7044, 
    7047, 
    7050, 
    7053, 
    7056, 
    7059, 
    7062, 
    7065, 
    7068, 
    7071, 
    7074, 
    7077, 
    7080, 
    7083, 
    7086, 
    7089, 
    7092, 
    7095, 
    7098, 
    7101, 
    7104, 
    7107, 
    7110, 
    7113, 
    7116, 
    7119, 
    7122, 
    7125, 
    7128, 
    7131, 
    7134, 
    7137, 
    7140, 
    7143, 
    7146, 
    7149, 
    7152, 
    7155, 
    7158, 
    7161, 
    7164, 
    7167, 
    7170, 
    7173, 
    7176, 
    7179, 
    7182, 
    7185, 
    7188, 
    7191, 
    7194, 
    7197, 
    7200, 
    7203, 
    7206, 
    7209, 
    7212, 
    7215, 
    7218, 
    7221, 
    7224, 
    7227, 
    7230, 
    7233, 
    7236, 
    7239, 
    7242, 
    7245, 
    7248, 
    7251, 
    7254, 
    7257, 
    7260, 
    7263, 
    7266, 
    7269, 
    7272, 
    7275, 
    7278, 
    7281, 
    7284, 
    7287, 
    7290, 
    7293, 
    7296, 
    7299, 
    7302, 
    7305, 
    7308, 
    7311, 
    7314, 
    7317, 
    7320, 
    7323, 
    7326, 
    7329, 
    7332, 
    7335, 
    7338, 
    7341, 
    7344, 
    7347, 
    7350, 
    7353, 
    7356, 
    7359, 
    7362, 
    7365, 
    7368, 
    7371, 
    7374, 
    7377, 
    7380, 
    7383, 
    7386, 
    7389, 
    7392, 
    7395, 
    7398, 
    7401, 
    7404, 
    7407, 
    7410, 
    7413, 
    7416, 
    7419, 
    7422, 
    7425, 
    7428, 
    7431, 
    7434, 
    7437, 
    7440, 
    7443, 
    7446, 
    7449, 
    7452, 
    7455, 
    7458, 
    7461, 
    7464, 
    7467, 
    7470, 
    7473, 
    7476, 
    7479, 
    7482, 
    7485, 
    7488, 
    7491, 
    7494, 
    7497, 
    7500, 
    7503, 
    7506, 
    7509, 
    7512, 
    7515, 
    7518, 
    7521, 
    7524, 
    7527, 
    7530, 
    7533, 
    7536, 
    7539, 
    7542, 
    7545, 
    7548, 
    7551, 
    7554, 
    7557, 
    7560, 
    7563, 
    7566, 
    7569, 
    7572, 
    7575, 
    7578, 
    7581, 
    7584, 
    7587, 
    7590, 
    7593, 
    7596, 
    7599, 
    7602, 
    7605, 
    7608, 
    7611, 
    7614, 
    7617, 
    7620, 
    7623, 
    7626, 
    7629, 
    7632, 
    7635, 
    7638, 
    7641, 
    7644, 
    7647, 
    7650, 
    7653, 
    7656, 
    7659, 
    7662, 
    7665, 
    7668, 
    7671, 
    7674, 
    7677, 
    7680, 
    7683, 
    7686, 
    7689, 
    7692, 
    7695, 
    7698, 
    7701, 
    7704, 
    7707, 
    7710, 
    7713, 
    7716, 
    7719, 
    7722, 
    7725, 
    7728, 
    7731, 
    7734, 
    7737, 
    7740, 
    7743, 
    7746, 
    7749, 
    7752, 
    7755, 
    7758, 
    7761, 
    7764, 
    7767, 
    7770, 
    7773, 
    7776, 
    7779, 
    7782, 
    7785, 
    7788, 
    7791, 
    7794, 
    7797, 
    7800, 
    7803, 
    7806, 
    7809, 
    7812, 
    7815, 
    7818, 
    7821, 
    7824, 
    7827, 
    7830, 
    7833, 
    7836, 
    7839, 
    7842, 
    7845, 
    7848, 
    7851, 
    7854, 
    7857, 
    7860, 
    7863, 
    7866, 
    7869, 
    7872, 
    7875, 
    7878, 
    7881, 
    7884, 
    7887, 
    7890, 
    7893, 
    7896, 
    7899, 
    7902, 
    7905, 
    7908, 
    7911, 
    7914, 
    7917, 
    7920, 
    7923, 
    7926, 
    7929, 
    7932, 
    7935, 
    7938, 
    7941, 
    7944, 
    7947, 
    7950, 
    7953, 
    7956, 
    7959, 
    7962, 
    7965, 
    7968, 
    7971, 
    7974, 
    7977, 
    7980, 
    7983, 
    7986, 
    7989, 
    7992, 
    7995, 
    7998, 
    8001, 
    8004, 
    8007, 
    8010, 
    8013, 
    8016, 
    8019, 
    8022, 
    8025, 
    8028, 
    8031, 
    8034, 
    8037, 
    8040, 
    8043, 
    8046, 
    8049, 
    8052, 
    8055, 
    8058, 
    8061, 
    8064, 
    8067, 
    8070, 
    8073, 
    8076, 
    8079, 
    8082, 
    8085, 
    8088, 
    8091, 
    8094, 
    8097, 
    8100, 
    8103, 
    8106, 
    8109, 
    8112, 
    8115, 
    8118, 
    8121, 
    8124, 
    8127, 
    8130, 
    8133, 
    8136, 
    8139, 
    8142, 
    8145, 
    8148, 
    8151, 
    8154, 
    8157, 
    8160, 
    8163, 
    8166, 
    8169, 
    8172, 
    8175, 
    8178, 
    8181, 
    8184, 
    8187, 
    8190, 
    8193, 
    8196, 
    8199, 
    8202, 
    8205, 
    8208, 
    8211, 
    8214, 
    8217, 
    8220, 
    8223, 
    8226, 
    8229, 
    8232, 
    8235, 
    8238, 
    8241, 
    8244, 
    8247, 
    8250, 
    8253, 
    8256, 
    8259, 
    8262, 
    8265, 
    8268, 
    8271, 
    8274, 
    8277, 
    8280, 
    8283, 
    8286, 
    8289, 
    8292, 
    8295, 
    8298, 
    8301, 
    8304, 
    8307, 
    8310, 
    8313, 
    8316, 
    8319, 
    8322, 
    8325, 
    8328, 
    8331, 
    8334, 
    8337, 
    8340, 
    8343, 
    8346, 
    8349, 
    8352, 
    8355, 
    8358, 
    8361, 
    8364, 
    8367, 
    8370, 
    8373, 
    8376, 
    8379, 
    8382, 
    8385, 
    8388, 
    8391, 
    8394, 
    8397, 
    8400, 
    8403, 
    8406, 
    8409, 
    8412, 
    8415, 
    8418, 
    8421, 
    8424, 
    8427, 
    8430, 
    8433, 
    8436, 
    8439, 
    8442, 
    8445, 
    8448, 
    8451, 
    8454, 
    8457, 
    8460, 
    8463, 
    8466, 
    8469, 
    8472, 
    8475, 
    8478, 
    8481, 
    8484, 
    8487, 
    8490, 
    8493, 
    8496, 
    8499, 
    8502, 
    8505, 
    8508, 
    8511, 
    8514, 
    8517, 
    8520, 
    8523, 
    8526, 
    8529, 
    8532, 
    8535, 
    8538, 
    8541, 
    8544, 
    8547, 
    8550, 
    8553, 
    8556, 
    8559, 
    8562, 
    8565, 
    8568, 
    8571, 
    8574, 
    8577, 
    8580, 
    8583, 
    8586, 
    8589, 
    8592, 
    8595, 
    8598, 
    8601, 
    8604, 
    8607, 
    8610, 
    8613, 
    8616, 
    8619, 
    8622, 
    8625, 
    8628, 
    8631, 
    8634, 
    8637, 
    8640, 
    8643, 
    8646, 
    8649, 
    8652, 
    8655, 
    8658, 
    8661, 
    8664, 
    8667, 
    8670, 
    8673, 
    8676, 
    8679, 
    8682, 
    8685, 
    8688, 
    8691, 
    8694, 
    8697, 
    8700, 
    8703, 
    8706, 
    8709, 
    8712, 
    8715, 
    8718, 
    8721, 
    8724, 
    8727, 
    8730, 
    8733, 
    8736, 
    8739, 
    8742, 
    8745, 
    8748, 
    8751, 
    8754, 
    8757, 
    8760, 
    8763, 
    8766, 
    8769, 
    8772, 
    8775, 
    8778, 
    8781, 
    8784, 
    8787, 
    8790, 
    8793, 
    8796, 
    8799, 
    8802, 
    8805, 
    8808, 
    8811, 
    8814, 
    8817, 
    8820, 
    8823, 
    8826, 
    8829, 
    8832, 
    8835, 
    8838, 
    8841, 
    8844, 
    8847, 
    8850, 
    8853, 
    8856, 
    8859, 
    8862, 
    8865, 
    8868, 
    8871, 
    8874, 
    8877, 
    8880, 
    8883, 
    8886, 
    8889, 
    8892, 
    8895, 
    8898, 
    8901, 
    8904, 
    8907, 
    8910, 
    8913, 
    8916, 
    8919, 
    8922, 
    8925, 
    8928, 
    8931, 
    8934, 
    8937, 
    8940, 
    8943, 
    8946, 
    8949, 
    8952, 
    8955, 
    8958, 
    8961, 
    8964, 
    8967, 
    8970, 
    8973, 
    8976, 
    8979, 
    8982, 
    8985, 
    8988, 
    8991, 
    8994, 
    8997, 
    9000, 
    9003, 
    9006, 
    9009, 
    9012, 
    9015, 
    9018, 
    9021, 
    9024, 
    9027, 
    9030, 
    9033, 
    9036, 
    9039, 
    9042, 
    9045, 
    9048, 
    9051, 
    9054, 
    9057, 
    9060, 
    9063, 
    9066, 
    9069, 
    9072, 
    9075, 
    9078, 
    9081, 
    9084, 
    9087, 
    9090, 
    9093, 
    9096, 
    9099, 
    9102, 
    9105, 
    9108, 
    9111, 
    9114, 
    9117, 
    9120, 
    9123, 
    9126, 
    9129, 
    9132, 
    9135, 
    9138, 
    9141, 
    9144, 
    9147, 
    9150, 
    9153, 
    9156, 
    9159, 
    9162, 
    9165, 
    9168, 
    9171, 
    9174, 
    9177, 
    9180, 
    9183, 
    9186, 
    9189, 
    9192, 
    9195, 
    9198, 
    9201, 
    9204, 
    9207, 
    9210, 
    9213, 
    9216, 
    9219, 
    9222, 
    9225, 
    9228, 
    9231, 
    9234, 
    9237, 
    9240, 
    9243, 
    9246, 
    9249, 
    9252, 
    9255, 
    9258, 
    9261, 
    9264, 
    9267, 
    9270, 
    9273, 
    9276, 
    9279, 
    9282, 
    9285, 
    9288, 
    9291, 
    9294, 
    9297, 
    9300, 
    9303, 
    9306, 
    9309, 
    9312, 
    9315, 
    9318, 
    9321, 
    9324, 
    9327, 
    9330, 
    9333, 
    9336, 
    9339, 
    9342, 
    9345, 
    9348, 
    9351, 
    9354, 
    9357, 
    9360, 
    9363, 
    9366, 
    9369, 
    9372, 
    9375, 
    9378, 
    9381, 
    9384, 
    9387, 
    9390, 
    9393, 
    9396, 
    9399, 
    9402, 
    9405, 
    9408, 
    9411, 
    9414, 
    9417, 
    9420, 
    9423, 
    9426, 
    9429, 
    9432, 
    9435, 
    9438, 
    9441, 
    9444, 
    9447, 
    9450, 
    9453, 
    9456, 
    9459, 
    9462, 
    9465, 
    9468, 
    9471, 
    9474, 
    9477, 
    9480, 
    9483, 
    9486, 
    9489, 
    9492, 
    9495, 
    9498, 
    9501, 
    9504, 
    9507, 
    9510, 
    9513, 
    9516, 
    9519, 
    9522, 
    9525, 
    9528, 
    9531, 
    9534, 
    9537, 
    9540, 
    9543, 
    9546, 
    9549, 
    9552, 
    9555, 
    9558, 
    9561, 
    9564, 
    9567, 
    9570, 
    9573, 
    9576, 
    9579, 
    9582, 
    9585, 
    9588, 
    9591, 
    9594, 
    9597, 
    9600, 
    9603, 
    9606, 
    9609, 
    9612, 
    9615, 
    9618, 
    9621, 
    9624, 
    9627, 
    9630, 
    9633, 
    9636, 
    9639, 
    9642, 
    9645, 
    9648, 
    9651, 
    9654, 
    9657, 
    9660, 
    9663, 
    9666, 
    9669, 
    9672, 
    9675, 
    9678, 
    9681, 
    9684, 
    9687, 
    9690, 
    9693, 
    9696, 
    9699, 
    9702, 
    9705, 
    9708, 
    9711, 
    9714, 
    9717, 
    9720, 
    9723, 
    9726, 
    9729, 
    9732, 
    9735, 
    9738, 
    9741, 
    9744, 
    9747, 
    9750, 
    9753, 
    9756, 
    9759, 
    9762, 
    9765, 
    9768, 
    9771, 
    9774, 
    9777, 
    9780, 
    9783, 
    9786, 
    9789, 
    9792, 
    9795, 
    9798, 
    9801, 
    9804, 
    9807, 
    9810, 
    9813, 
    9816, 
    9819, 
    9822, 
    9825, 
    9828, 
    9831, 
    9834, 
    9837, 
    9840, 
    9843, 
    9846, 
    9849, 
    9852, 
    9855, 
    9858, 
    9861, 
    9864, 
    9867, 
    9870, 
    9873, 
    9876, 
    9879, 
    9882, 
    9885, 
    9888, 
    9891, 
    9894, 
    9897, 
    9900, 
    9903, 
    9906, 
    9909, 
    9912, 
    9915, 
    9918, 
    9921, 
    9924, 
    9927, 
    9930, 
    9933, 
    9936, 
    9939, 
    9942, 
    9945, 
    9948, 
    9951, 
    9954, 
    9957, 
    9960, 
    9963, 
    9966, 
    9969, 
    9972, 
    9975, 
    9978, 
    9981, 
    9984, 
    9987, 
    9990, 
    9993, 
    9996, 
    9999, 
    10002, 
    10005, 
    10008, 
    10011, 
    10014, 
    10017, 
    10020, 
    10023, 
    10026, 
    10029, 
    10032, 
    10035, 
    10038, 
    10041, 
    10044, 
    10047, 
    10050, 
    10053, 
    10056, 
    10059, 
    10062, 
    10065, 
    10068, 
    10071, 
    10074, 
    10077, 
    10080, 
    10083, 
    10086, 
    10089, 
    10092, 
    10095, 
    10098, 
    10101, 
    10104, 
    10107, 
    10110, 
    10113, 
    10116, 
    10119, 
    10122, 
    10125, 
    10128, 
    10131, 
    10134, 
    10137, 
    10140, 
    10143, 
    10146, 
    10149, 
    10152, 
    10155, 
    10158, 
    10161, 
    10164, 
    10167, 
    10170, 
    10173, 
    10176, 
    10179, 
    10182, 
    10185, 
    10188, 
    10191, 
    10194, 
    10197, 
    10200, 
    10203, 
    10206, 
    10209, 
    10212, 
    10215, 
    10218, 
    10221, 
    10224, 
    10227, 
    10230, 
    10233, 
    10236, 
    10239, 
    10242, 
    10245, 
    10248, 
    10251, 
    10254, 
    10257, 
    10260, 
    10263, 
    10266, 
    10269, 
    10272, 
    10275, 
    10278, 
    10281, 
    10284, 
    10287, 
    10290, 
    10293, 
    10296, 
    10299, 
    10302, 
    10305, 
    10308, 
    10311, 
    10314, 
    10317, 
    10320, 
    10323, 
    10326, 
    10329, 
    10332, 
    10335, 
    10338, 
    10341, 
    10344, 
    10347, 
    10350, 
    10353, 
    10356, 
    10359, 
    10362, 
    10365, 
    10368, 
    10371, 
    10374, 
    10377, 
    10380, 
    10383, 
    10386, 
    10389, 
    10392, 
    10395, 
    10398, 
    10401, 
    10404, 
    10407, 
    10410, 
    10413, 
    10416, 
    10419, 
    10422, 
    10425, 
    10428, 
    10431, 
    10434, 
    10437, 
    10440, 
    10443, 
    10446, 
    10449, 
    10452, 
    10455, 
    10458, 
    10461, 
    10464, 
    10467, 
    10470, 
    10473, 
    10476, 
    10479, 
    10482, 
    10485, 
    10488, 
    10491, 
    10494, 
    10497, 
    10500, 
    10503, 
    10506, 
    10509, 
    10512, 
    10515, 
    10518, 
    10521, 
    10524, 
    10527, 
    10530, 
    10533, 
    10536, 
    10539, 
    10542, 
    10545, 
    10548, 
    10551, 
    10554, 
    10557, 
    10560, 
    10563, 
    10566, 
    10569, 
    10572, 
    10575, 
    10578, 
    10581, 
    10584, 
    10587, 
    10590, 
    10593, 
    10596, 
    10599, 
    10602, 
    10605, 
    10608, 
    10611, 
    10614, 
    10617, 
    10620, 
    10623, 
    10626, 
    10629, 
    10632, 
    10635, 
    10638, 
    10641, 
    10644, 
    10647, 
    10650, 
    10653, 
    10656, 
    10659, 
    10662, 
    10665, 
    10668, 
    10671, 
    10674, 
    10677, 
    10680, 
    10683, 
    10686, 
    10689, 
    10692, 
    10695, 
    10698, 
    10701, 
    10704, 
    10707, 
    10710, 
    10713, 
    10716, 
    10719, 
    10722, 
    10725, 
    10728, 
    10731, 
    10734, 
    10737, 
    10740, 
    10743, 
    10746, 
    10749, 
    10752, 
    10755, 
    10758, 
    10761, 
    10764, 
    10767, 
    10770, 
    10773, 
    10776, 
    10779, 
    10782, 
    10785, 
    10788, 
    10791, 
    10794, 
    10797, 
    10800, 
    10803, 
    10806, 
    10809, 
    10812, 
    10815, 
    10818, 
    10821, 
    10824, 
    10827, 
    10830, 
    10833, 
    10836, 
    10839, 
    10842, 
    10845, 
    10848, 
    10851, 
    10854, 
    10857, 
    10860, 
    10863, 
    10866, 
    10869, 
    10872, 
    10875, 
    10878, 
    10881, 
    10884, 
    10887, 
    10890, 
    10893, 
    10896, 
    10899, 
    10902, 
    10905, 
    10908, 
    10911, 
    10914, 
    10917, 
    10920, 
    10923, 
    10926, 
    10929, 
    10932, 
    10935, 
    10938, 
    10941, 
    10944, 
    10947, 
    10950, 
    10953, 
    10956, 
    10959, 
    10962, 
    10965, 
    10968, 
    10971, 
    10974, 
    10977, 
    10980, 
    10983, 
    10986, 
    10989, 
    10992, 
    10995, 
    10998, 
    11001, 
    11004, 
    11007, 
    11010, 
    11013, 
    11016, 
    11019, 
    11022, 
    11025, 
    11028, 
    11031, 
    11034, 
    11037, 
    11040, 
    11043, 
    11046, 
    11049, 
    11052, 
    11055, 
    11058, 
    11061, 
    11064, 
    11067, 
    11070, 
    11073, 
    11076, 
    11079, 
    11082, 
    11085, 
    11088, 
    11091, 
    11094, 
    11097, 
    11100, 
    11103, 
    11106, 
    11109, 
    11112, 
    11115, 
    11118, 
    11121, 
    11124, 
    11127, 
    11130, 
    11133, 
    11136, 
    11139, 
    11142, 
    11145, 
    11148, 
    11151, 
    11154, 
    11157, 
    11160, 
    11163, 
    11166, 
    11169, 
    11172, 
    11175, 
    11178, 
    11181, 
    11184, 
    11187, 
    11190, 
    11193, 
    11196, 
    11199, 
    11202, 
    11205, 
    11208, 
    11211, 
    11214, 
    11217, 
    11220, 
    11223, 
    11226, 
    11229, 
    11232, 
    11235, 
    11238, 
    11241, 
    11244, 
    11247, 
    11250, 
    11253, 
    11256, 
    11259, 
    11262, 
    11265, 
    11268, 
    11271, 
    11274, 
    11277, 
    11280, 
    11283, 
    11286, 
    11289, 
    11292, 
    11295, 
    11298, 
    11301, 
    11304, 
    11307, 
    11310, 
    11313, 
    11316, 
    11319, 
    11322, 
    11325, 
    11328, 
    11331, 
    11334, 
    11337, 
    11340, 
    11343, 
    11346, 
    11349, 
    11352, 
    11355, 
    11358, 
    11361, 
    11364, 
    11367, 
    11370, 
    11373, 
    11376, 
    11379, 
    11382, 
    11385, 
    11388, 
    11391, 
    11394, 
    11397, 
    11400, 
    11403, 
    11406, 
    11409, 
    11412, 
    11415, 
    11418, 
    11421, 
    11424, 
    11427, 
    11430, 
    11433, 
    11436, 
    11439, 
    11442, 
    11445, 
    11448, 
    11451, 
    11454, 
    11457, 
    11460, 
    11463, 
    11466, 
    11469, 
    11472, 
    11475, 
    11478, 
    11481, 
    11484, 
    11487, 
    11490, 
    11493, 
    11496, 
    11499, 
    11502, 
    11505, 
    11508, 
    11511, 
    11514, 
    11517, 
    11520, 
    11523, 
    11526, 
    11529, 
    11532, 
    11535, 
    11538, 
    11541, 
    11544, 
    11547, 
    11550, 
    11553, 
    11556, 
    11559, 
    11562, 
    11565, 
    11568, 
    11571, 
    11574, 
    11577, 
    11580, 
    11583, 
    11586, 
    11589, 
    11592, 
    11595, 
    11598, 
    11601, 
    11604, 
    11607, 
    11610, 
    11613, 
    11616, 
    11619, 
    11622, 
    11625, 
    11628, 
    11631, 
    11634, 
    11637, 
    11640, 
    11643, 
    11646, 
    11649, 
    11652, 
    11655, 
    11658, 
    11661, 
    11664, 
    11667, 
    11670, 
    11673, 
    11676, 
    11679, 
    11682, 
    11685, 
    11688, 
    11691, 
    11694, 
    11697, 
    11700, 
    11703, 
    11706, 
    11709, 
    11712, 
    11715, 
    11718, 
    11721, 
    11724, 
    11727, 
    11730, 
    11733, 
    11736, 
    11739, 
    11742, 
    11745, 
    11748, 
    11751, 
    11754, 
    11757, 
    11760, 
    11763, 
    11766, 
    11769, 
    11772, 
    11775, 
    11778, 
    11781, 
    11784, 
    11787, 
    11790, 
    11793, 
    11796, 
    11799, 
    11802, 
    11805, 
    11808, 
    11811, 
    11814, 
    11817, 
    11820, 
    11823, 
    11826, 
    11829, 
    11832, 
    11835, 
    11838, 
    11841, 
    11844, 
    11847, 
    11850, 
    11853, 
    11856, 
    11859, 
    11862, 
    11865, 
    11868, 
    11871, 
    11874, 
    11877, 
    11880, 
    11883, 
    11886, 
    11889, 
    11892, 
    11895, 
    11898, 
    11901, 
    11904, 
    11907, 
    11910, 
    11913, 
    11916, 
    11919, 
    11922, 
    11925, 
    11928, 
    11931, 
    11934, 
    11937, 
    11940, 
    11943, 
    11946, 
    11949, 
    11952, 
    11955, 
    11958, 
    11961, 
    11964, 
    11967, 
    11970, 
    11973, 
    11976, 
    11979, 
    11982, 
    11985, 
    11988, 
    11991, 
    11994, 
    11997, 
    12000, 
    12003, 
    12006, 
    12009, 
    12012, 
    12015, 
    12018, 
    12021, 
    12024, 
    12027, 
    12030, 
    12033, 
    12036, 
    12039, 
    12042, 
    12045, 
    12048, 
    12051, 
    12054, 
    12057, 
    12060, 
    12063, 
    12066, 
    12069, 
    12072, 
    12075, 
    12078, 
    12081, 
    12084, 
    12087, 
    12090, 
    12093, 
    12096, 
    12099, 
    12102, 
    12105, 
    12108, 
    12111, 
    12114, 
    12117, 
    12120, 
    12123, 
    12126, 
    12129, 
    12132, 
    12135, 
    12138, 
    12141, 
    12144, 
    12147, 
    12150, 
    12153, 
    12156, 
    12159, 
    12162, 
    12165, 
    12168, 
    12171, 
    12174, 
    12177, 
    12180, 
    12183, 
    12186, 
    12189, 
    12192, 
    12195, 
    12198, 
    12201, 
    12204, 
    12207, 
    12210, 
    12213, 
    12216, 
    12219, 
    12222, 
    12225, 
    12228, 
    12231, 
    12234, 
    12237, 
    12240, 
    12243, 
    12246, 
    12249, 
    12252, 
    12255, 
    12258, 
    12261, 
    12264, 
    12267, 
    12270, 
    12273, 
    12276, 
    12279, 
    12282, 
    12285, 
    12288, 
    12291, 
    12294, 
    12297, 
    12300, 
    12303, 
    12306, 
    12309, 
    12312, 
    12315, 
    12318, 
    12321, 
    12324, 
    12327, 
    12330, 
    12333, 
    12336, 
    12339, 
    12342, 
    12345, 
    12348, 
    12351, 
    12354, 
    12357, 
    12360, 
    12363, 
    12366, 
    12369, 
    12372, 
    12375, 
    12378, 
    12381, 
    12384, 
    12387, 
    12390, 
    12393, 
    12396, 
    12399, 
    12402, 
    12405, 
    12408, 
    12411, 
    12414, 
    12417, 
    12420, 
    12423, 
    12426, 
    12429, 
    12432, 
    12435, 
    12438, 
    12441, 
    12444, 
    12447, 
    12450, 
    12453, 
    12456, 
    12459, 
    12462, 
    12465, 
    12468, 
    12471, 
    12474, 
    12477, 
    12480, 
    12483, 
    12486, 
    12489, 
    12492, 
    12495, 
    12498, 
    12501, 
    12504, 
    12507, 
    12510, 
    12513, 
    12516, 
    12519, 
    12522, 
    12525, 
    12528, 
    12531, 
    12534, 
    12537, 
    12540, 
    12543, 
    12546, 
    12549, 
    12552, 
    12555, 
    12558, 
    12561, 
    12564, 
    12567, 
    12570, 
    12573, 
    12576, 
    12579, 
    12582, 
    12585, 
    12588, 
    12591, 
    12594, 
    12597, 
    12600, 
    12603, 
    12606, 
    12609, 
    12612, 
    12615, 
    12618, 
    12621, 
    12624, 
    12627, 
    12630, 
    12633, 
    12636, 
    12639, 
    12642, 
    12645, 
    12648, 
    12651, 
    12654, 
    12657, 
    12660, 
    12663, 
    12666, 
    12669, 
    12672, 
    12675, 
    12678, 
    12681, 
    12684, 
    12687, 
    12690, 
    12693, 
    12696, 
    12699, 
    12702, 
    12705, 
    12708, 
    12711, 
    12714, 
    12717, 
    12720, 
    12723, 
    12726, 
    12729, 
    12732, 
    12735, 
    12738, 
    12741, 
    12744, 
    12747, 
    12750, 
    12753, 
    12756, 
    12759, 
    12762, 
    12765, 
    12768, 
    12771, 
    12774, 
    12777, 
    12780, 
    12783, 
    12786, 
    12789, 
    12792, 
    12795, 
    12798, 
    12801, 
    12804, 
    12807, 
    12810, 
    12813, 
    12816, 
    12819, 
    12822, 
    12825, 
    12828, 
    12831, 
    12834, 
    12837, 
    12840, 
    12843, 
    12846, 
    12849, 
    12852, 
    12855, 
    12858, 
    12861, 
    12864, 
    12867, 
    12870, 
    12873, 
    12876, 
    12879, 
    12882, 
    12885, 
    12888, 
    12891, 
    12894, 
    12897, 
    12900, 
    12903, 
    12906, 
    12909, 
    12912, 
    12915, 
    12918, 
    12921, 
    12924, 
    12927, 
    12930, 
    12933, 
    12936, 
    12939, 
    12942, 
    12945, 
    12948, 
    12951, 
    12954, 
    12957, 
    12960, 
    12963, 
    12966, 
    12969, 
    12972, 
    12975, 
    12978, 
    12981, 
    12984, 
    12987, 
    12990, 
    12993, 
    12996, 
    12999, 
    13002, 
    13005, 
    13008, 
    13011, 
    13014, 
    13017, 
    13020, 
    13023, 
    13026, 
    13029, 
    13032, 
    13035, 
    13038, 
    13041, 
    13044, 
    13047, 
    13050, 
    13053, 
    13056, 
    13059, 
    13062, 
    13065, 
    13068, 
    13071, 
    13074, 
    13077, 
    13080, 
    13083, 
    13086, 
    13089, 
    13092, 
    13095, 
    13098, 
    13101, 
    13104, 
    13107, 
    13110, 
    13113, 
    13116, 
    13119, 
    13122, 
    13125, 
    13128, 
    13131, 
    13134, 
    13137, 
    13140, 
    13143, 
    13146, 
    13149, 
    13152, 
    13155, 
    13158, 
    13161, 
    13164, 
    13167, 
    13170, 
    13173, 
    13176, 
    13179, 
    13182, 
    13185, 
    13188, 
    13191, 
    13194, 
    13197, 
    13200, 
    13203, 
    13206, 
    13209, 
    13212, 
    13215, 
    13218, 
    13221, 
    13224, 
    13227, 
    13230, 
    13233, 
    13236, 
    13239, 
    13242, 
    13245, 
    13248, 
    13251, 
    13254, 
    13257, 
    13260, 
    13263, 
    13266, 
    13269, 
    13272, 
    13275, 
    13278, 
    13281, 
    13284, 
    13287, 
    13290, 
    13293, 
    13296, 
    13299, 
    13302, 
    13305, 
    13308, 
    13311, 
    13314, 
    13317, 
    13320, 
    13323, 
    13326, 
    13329, 
    13332, 
    13335, 
    13338, 
    13341, 
    13344, 
    13347, 
    13350, 
    13353, 
    13356, 
    13359, 
    13362, 
    13365, 
    13368, 
    13371, 
    13374, 
    13377, 
    13380, 
    13383, 
    13386, 
    13389, 
    13392, 
    13395, 
    13398, 
    13401, 
    13404, 
    13407, 
    13410, 
    13413, 
    13416, 
    13419, 
    13422, 
    13425, 
    13428, 
    13431, 
    13434, 
    13437, 
    13440, 
    13443, 
    13446, 
    13449, 
    13452, 
    13455, 
    13458, 
    13461, 
    13464, 
    13467, 
    13470, 
    13473, 
    13476, 
    13479, 
    13482, 
    13485, 
    13488, 
    13491, 
    13494, 
    13497, 
    13500, 
    13503, 
    13506, 
    13509, 
    13512, 
    13515, 
    13518, 
    13521, 
    13524, 
    13527, 
    13530, 
    13533, 
    13536, 
    13539, 
    13542, 
    13545, 
    13548, 
    13551, 
    13554, 
    13557, 
    13560, 
    13563, 
    13566, 
    13569, 
    13572, 
    13575, 
    13578, 
    13581, 
    13584, 
    13587, 
    13590, 
    13593, 
    13596, 
    13599, 
    13602, 
    13605, 
    13608, 
    13611, 
    13614, 
    13617, 
    13620, 
    13623, 
    13626, 
    13629, 
    13632, 
    13635, 
    13638, 
    13641, 
    13644, 
    13647, 
    13650, 
    13653, 
    13656, 
    13659, 
    13662, 
    13665, 
    13668, 
    13671, 
    13674, 
    13677, 
    13680, 
    13683, 
    13686, 
    13689, 
    13692, 
    13695, 
    13698, 
    13701, 
    13704, 
    13707, 
    13710, 
    13713, 
    13716, 
    13719, 
    13722, 
    13725, 
    13728, 
    13731, 
    13734, 
    13737, 
    13740, 
    13743, 
    13746, 
    13749, 
    13752, 
    13755, 
    13758, 
    13761, 
    13764, 
    13767, 
    13770, 
    13773, 
    13776, 
    13779, 
    13782, 
    13785, 
    13788, 
    13791, 
    13794, 
    13797, 
    13800, 
    13803, 
    13806, 
    13809, 
    13812, 
    13815, 
    13818, 
    13821, 
    13824, 
    13827, 
    13830, 
    13833, 
    13836, 
    13839, 
    13842, 
    13845, 
    13848, 
    13851, 
    13854, 
    13857, 
    13860, 
    13863, 
    13866, 
    13869, 
    13872, 
    13875, 
    13878, 
    13881, 
    13884, 
    13887, 
    13890, 
    13893, 
    13896, 
    13899, 
    13902, 
    13905, 
    13908, 
    13911, 
    13914, 
    13917, 
    13920, 
    13923, 
    13926, 
    13929, 
    13932, 
    13935, 
    13938, 
    13941, 
    13944, 
    13947, 
    13950, 
    13953, 
    13956, 
    13959, 
    13962, 
    13965, 
    13968, 
    13971, 
    13974, 
    13977, 
    13980, 
    13983, 
    13986, 
    13989, 
    13992, 
    13995, 
    13998, 
    14001, 
    14004, 
    14007, 
    14010, 
    14013, 
    14016, 
    14019, 
    14022, 
    14025, 
    14028, 
    14031, 
    14034, 
    14037, 
    14040, 
    14043, 
    14046, 
    14049, 
    14052, 
    14055, 
    14058, 
    14061, 
    14064, 
    14067, 
    14070, 
    14073, 
    14076, 
    14079, 
    14082, 
    14085, 
    14088, 
    14091, 
    14094, 
    14097, 
    14100, 
    14103, 
    14106, 
    14109, 
    14112, 
    14115, 
    14118, 
    14121, 
    14124, 
    14127, 
    14130, 
    14133, 
    14136, 
    14139, 
    14142, 
    14145, 
    14148, 
    14151, 
    14154, 
    14157, 
    14160, 
    14163, 
    14166, 
    14169, 
    14172, 
    14175, 
    14178, 
    14181, 
    14184, 
    14187, 
    14190, 
    14193, 
    14196, 
    14199, 
    14202, 
    14205, 
    14208, 
    14211, 
    14214, 
    14217, 
    14220, 
    14223, 
    14226, 
    14229, 
    14232, 
    14235, 
    14238, 
    14241, 
    14244, 
    14247, 
    14250, 
    14253, 
    14256, 
    14259, 
    14262, 
    14265, 
    14268, 
    14271, 
    14274, 
    14277, 
    14280, 
    14283, 
    14286, 
    14289, 
    14292, 
    14295, 
    14298, 
    14301, 
    14304, 
    14307, 
    14310, 
    14313, 
    14316, 
    14319, 
    14322, 
    14325, 
    14328, 
    14331, 
    14334, 
    14337, 
    14340, 
    14343, 
    14346, 
    14349, 
    14352, 
    14355, 
    14358, 
    14361, 
    14364, 
    14367, 
    14370, 
    14373, 
    14376, 
    14379, 
    14382, 
    14385, 
    14388, 
    14391, 
    14394, 
    14397, 
    14400, 
    14403, 
    14406, 
    14409, 
    14412, 
    14415, 
    14418, 
    14421, 
    14424, 
    14427, 
    14430, 
    14433, 
    14436, 
    14439, 
    14442, 
    14445, 
    14448, 
    14451, 
    14454, 
    14457, 
    14460, 
    14463, 
    14466, 
    14469, 
    14472, 
    14475, 
    14478, 
    14481, 
    14484, 
    14487, 
    14490, 
    14493, 
    14496, 
    14499, 
    14502, 
    14505, 
    14508, 
    14511, 
    14514, 
    14517, 
    14520, 
    14523, 
    14526, 
    14529, 
    14532, 
    14535, 
    14538, 
    14541, 
    14544, 
    14547, 
    14550, 
    14553, 
    14556, 
    14559, 
    14562, 
    14565, 
    14568, 
    14571, 
    14574, 
    14577, 
    14580, 
    14583, 
    14586, 
    14589, 
    14592, 
    14595, 
    14598, 
    14601, 
    14604, 
    14607, 
    14610, 
    14613, 
    14616, 
    14619, 
    14622, 
    14625, 
    14628, 
    14631, 
    14634, 
    14637, 
    14640, 
    14643, 
    14646, 
    14649, 
    14652, 
    14655, 
    14658, 
    14661, 
    14664, 
    14667, 
    14670, 
    14673, 
    14676, 
    14679, 
    14682, 
    14685, 
    14688, 
    14691, 
    14694, 
    14697, 
    14700, 
    14703, 
    14706, 
    14709, 
    14712, 
    14715, 
    14718, 
    14721, 
    14724, 
    14727, 
    14730, 
    14733, 
    14736, 
    14739, 
    14742, 
    14745, 
    14748, 
    14751, 
    14754, 
    14757, 
    14760, 
    14763, 
    14766, 
    14769, 
    14772, 
    14775, 
    14778, 
    14781, 
    14784, 
    14787, 
    14790, 
    14793, 
    14796, 
    14799, 
    14802, 
    14805, 
    14808, 
    14811, 
    14814, 
    14817, 
    14820, 
    14823, 
    14826, 
    14829, 
    14832, 
    14835, 
    14838, 
    14841, 
    14844, 
    14847, 
    14850, 
    14853, 
    14856, 
    14859, 
    14862, 
    14865, 
    14868, 
    14871, 
    14874, 
    14877, 
    14880, 
    14883, 
    14886, 
    14889, 
    14892, 
    14895, 
    14898, 
    14901, 
    14904, 
    14907, 
    14910, 
    14913, 
    14916, 
    14919, 
    14922, 
    14925, 
    14928, 
    14931, 
    14934, 
    14937, 
    14940, 
    14943, 
    14946, 
    14949, 
    14952, 
    14955, 
    14958, 
    14961, 
    14964, 
    14967, 
    14970, 
    14973, 
    14976, 
    14979, 
    14982, 
    14985, 
    14988, 
    14991, 
    14994, 
    14997, 
    15000, 
    15003, 
    15006, 
    15009, 
    15012, 
    15015, 
    15018, 
    15021, 
    15024, 
    15027, 
    15030, 
    15033, 
    15036, 
    15039, 
    15042, 
    15045, 
    15048, 
    15051, 
    15054, 
    15057, 
    15060, 
    15063, 
    15066, 
    15069, 
    15072, 
    15075, 
    15078, 
    15081, 
    15084, 
    15087, 
    15090, 
    15093, 
    15096, 
    15099, 
    15102, 
    15105, 
    15108, 
    15111, 
    15114, 
    15117, 
    15120, 
    15123, 
    15126, 
    15129, 
    15132, 
    15135, 
    15138, 
    15141, 
    15144, 
    15147, 
    15150, 
    15153, 
    15156, 
    15159, 
    15162, 
    15165, 
    15168, 
    15171, 
    15174, 
    15177, 
    15180, 
    15183, 
    15186, 
    15189, 
    15192, 
    15195, 
    15198, 
    15201, 
    15204, 
    15207, 
    15210, 
    15213, 
    15216, 
    15219, 
    15222, 
    15225, 
    15228, 
    15231, 
    15234, 
    15237, 
    15240, 
    15243, 
    15246, 
    15249, 
    15252, 
    15255, 
    15258, 
    15261, 
    15264, 
    15267, 
    15270, 
    15273, 
    15276, 
    15279, 
    15282, 
    15285, 
    15288, 
    15291, 
    15294, 
    15297, 
    15300, 
    15303, 
    15306, 
    15309, 
    15312, 
    15315, 
    15318, 
    15321, 
    15324, 
    15327, 
    15330, 
    15333, 
    15336, 
    15339, 
    15342, 
    15345, 
    15348, 
    15351, 
    15354, 
    15357, 
    15360, 
    15363, 
    15366, 
    15369, 
    15372, 
    15375, 
    15378, 
    15381, 
    15384, 
    15387, 
    15390, 
    15393, 
    15396, 
    15399, 
    15402, 
    15405, 
    15408, 
    15411, 
    15414, 
    15417, 
    15420, 
    15423, 
    15426, 
    15429, 
    15432, 
    15435, 
    15438, 
    15441, 
    15444, 
    15447, 
    15450, 
    15453, 
    15456, 
    15459, 
    15462, 
    15465, 
    15468, 
    15471, 
    15474, 
    15477, 
    15480, 
    15483, 
    15486, 
    15489, 
    15492, 
    15495, 
    15498, 
    15501, 
    15504, 
    15507, 
    15510, 
    15513, 
    15516, 
    15519, 
    15522, 
    15525, 
    15528, 
    15531, 
    15534, 
    15537, 
    15540, 
    15543, 
    15546, 
    15549, 
    15552, 
    15555, 
    15558, 
    15561, 
    15564, 
    15567, 
    15570, 
    15573, 
    15576, 
    15579, 
    15582, 
    15585, 
    15588, 
    15591, 
    15594, 
    15597, 
    15600, 
    15603, 
    15606, 
    15609, 
    15612, 
    15615, 
    15618, 
    15621, 
    15624, 
    15627, 
    15630, 
    15633, 
    15636, 
    15639, 
    15642, 
    15645, 
    15648, 
    15651, 
    15654, 
    15657, 
    15660, 
    15663, 
    15666, 
    15669, 
    15672, 
    15675, 
    15678, 
    15681, 
    15684, 
    15687, 
    15690, 
    15693, 
    15696, 
    15699, 
    15702, 
    15705, 
    15708, 
    15711, 
    15714, 
    15717, 
    15720, 
    15723, 
    15726, 
    15729, 
    15732, 
    15735, 
    15738, 
    15741, 
    15744, 
    15747, 
    15750, 
    15753, 
    15756, 
    15759, 
    15762, 
    15765, 
    15768, 
    15771, 
    15774, 
    15777, 
    15780, 
    15783, 
    15786, 
    15789, 
    15792, 
    15795, 
    15798, 
    15801, 
    15804, 
    15807, 
    15810, 
    15813, 
    15816, 
    15819, 
    15822, 
    15825, 
    15828, 
    15831, 
    15834, 
    15837, 
    15840, 
    15843, 
    15846, 
    15849, 
    15852, 
    15855, 
    15858, 
    15861, 
    15864, 
    15867, 
    15870, 
    15873, 
    15876, 
    15879, 
    15882, 
    15885, 
    15888, 
    15891, 
    15894, 
    15897, 
    15900, 
    15903, 
    15906, 
    15909, 
    15912, 
    15915, 
    15918, 
    15921, 
    15924, 
    15927, 
    15930, 
    15933, 
    15936, 
    15939, 
    15942, 
    15945, 
    15948, 
    15951, 
    15954, 
    15957, 
    15960, 
    15963, 
    15966, 
    15969, 
    15972, 
    15975, 
    15978, 
    15981, 
    15984, 
    15987, 
    15990, 
    15993, 
    15996, 
    15999, 
    16002, 
    16005, 
    16008, 
    16011, 
    16014, 
    16017, 
    16020, 
    16023, 
    16026, 
    16029, 
    16032, 
    16035, 
    16038, 
    16041, 
    16044, 
    16047, 
    16050, 
    16053, 
    16056, 
    16059, 
    16062, 
    16065, 
    16068, 
    16071, 
    16074, 
    16077, 
    16080, 
    16083, 
    16086, 
    16089, 
    16092, 
    16095, 
    16098, 
    16101, 
    16104, 
    16107, 
    16110, 
    16113, 
    16116, 
    16119, 
    16122, 
    16125, 
    16128, 
    16131, 
    16134, 
    16137, 
    16140, 
    16143, 
    16146, 
    16149, 
    16152, 
    16155, 
    16158, 
    16161, 
    16164, 
    16167, 
    16170, 
    16173, 
    16176, 
    16179, 
    16182, 
    16185, 
    16188, 
    16191, 
    16194, 
    16197, 
    16200, 
    16203, 
    16206, 
    16209, 
    16212, 
    16215, 
    16218, 
    16221, 
    16224, 
    16227, 
    16230, 
    16233, 
    16236, 
    16239, 
    16242, 
    16245, 
    16248, 
    16251, 
    16254, 
    16257, 
    16260, 
    16263, 
    16266, 
    16269, 
    16272, 
    16275, 
    16278, 
    16281, 
    16284, 
    16287, 
    16290, 
    16293, 
    16296, 
    16299, 
    16302, 
    16305, 
    16308, 
    16311, 
    16314, 
    16317, 
    16320, 
    16323, 
    16326, 
    16329, 
    16332, 
    16335, 
    16338, 
    16341, 
    16344, 
    16347, 
    16350, 
    16353, 
    16356, 
    16359, 
    16362, 
    16365, 
    16368, 
    16371, 
    16374, 
    16377, 
    16380, 
    16383, 
    16386, 
    16389, 
    16392, 
    16395, 
    16398, 
    16401, 
    16404, 
    16407, 
    16410, 
    16413, 
    16416, 
    16419, 
    16422, 
    16425, 
    16428, 
    16431, 
    16434, 
    16437, 
    16440, 
    16443, 
    16446, 
    16449, 
    16452, 
    16455, 
    16458, 
    16461, 
    16464, 
    16467, 
    16470, 
    16473, 
    16476, 
    16479, 
    16482, 
    16485, 
    16488, 
    16491, 
    16494, 
    16497, 
    16500, 
    16503, 
    16506, 
    16509, 
    16512, 
    16515, 
    16518, 
    16521, 
    16524, 
    16527, 
    16530, 
    16533, 
    16536, 
    16539, 
    16542, 
    16545, 
    16548, 
    16551, 
    16554, 
    16557, 
    16560, 
    16563, 
    16566, 
    16569, 
    16572, 
    16575, 
    16578, 
    16581, 
    16584, 
    16587, 
    16590, 
    16593, 
    16596, 
    16599, 
    16602, 
    16605, 
    16608, 
    16611, 
    16614, 
    16617, 
    16620, 
    16623, 
    16626, 
    16629, 
    16632, 
    16635, 
    16638, 
    16641, 
    16644, 
    16647, 
    16650, 
    16653, 
    16656, 
    16659, 
    16662, 
    16665, 
    16668, 
    16671, 
    16674, 
    16677, 
    16680, 
    16683, 
    16686, 
    16689, 
    16692, 
    16695, 
    16698, 
    16701, 
    16704, 
    16707, 
    16710, 
    16713, 
    16716, 
    16719, 
    16722, 
    16725, 
    16728, 
    16731, 
    16734, 
    16737, 
    16740, 
    16743, 
    16746, 
    16749, 
    16752, 
    16755, 
    16758, 
    16761, 
    16764, 
    16767, 
    16770, 
    16773, 
    16776, 
    16779, 
    16782, 
    16785, 
    16788, 
    16791, 
    16794, 
    16797, 
    16800, 
    16803, 
    16806, 
    16809, 
    16812, 
    16815, 
    16818, 
    16821, 
    16824, 
    16827, 
    16830, 
    16833, 
    16836, 
    16839, 
    16842, 
    16845, 
    16848, 
    16851, 
    16854, 
    16857, 
    16860, 
    16863, 
    16866, 
    16869, 
    16872, 
    16875, 
    16878, 
    16881, 
    16884, 
    16887, 
    16890, 
    16893, 
    16896, 
    16899, 
    16902, 
    16905, 
    16908, 
    16911, 
    16914, 
    16917, 
    16920, 
    16923, 
    16926, 
    16929, 
    16932, 
    16935, 
    16938, 
    16941, 
    16944, 
    16947, 
    16950, 
    16953, 
    16956, 
    16959, 
    16962, 
    16965, 
    16968, 
    16971, 
    16974, 
    16977, 
    16980, 
    16983, 
    16986, 
    16989, 
    16992, 
    16995, 
    16998, 
    17001, 
    17004, 
    17007, 
    17010, 
    17013, 
    17016, 
    17019, 
    17022, 
    17025, 
    17028, 
    17031, 
    17034, 
    17037, 
    17040, 
    17043, 
    17046, 
    17049, 
    17052, 
    17055, 
    17058, 
    17061, 
    17064, 
    17067, 
    17070, 
    17073, 
    17076, 
    17079, 
    17082, 
    17085, 
    17088, 
    17091, 
    17094, 
    17097, 
    17100, 
    17103, 
    17106, 
    17109, 
    17112, 
    17115, 
    17118, 
    17121, 
    17124, 
    17127, 
    17130, 
    17133, 
    17136, 
    17139, 
    17142, 
    17145, 
    17148, 
    17151, 
    17154, 
    17157, 
    17160, 
    17163, 
    17166, 
    17169, 
    17172, 
    17175, 
    17178, 
    17181, 
    17184, 
    17187, 
    17190, 
    17193, 
    17196, 
    17199, 
    17202, 
    17205, 
    17208, 
    17211, 
    17214, 
    17217, 
    17220, 
    17223, 
    17226, 
    17229, 
    17232, 
    17235, 
    17238, 
    17241, 
    17244, 
    17247, 
    17250, 
    17253, 
    17256, 
    17259, 
    17262, 
    17265, 
    17268, 
    17271, 
    17274, 
    17277, 
    17280, 
    17283, 
    17286, 
    17289, 
    17292, 
    17295, 
    17298, 
    17301, 
    17304, 
    17307, 
    17310, 
    17313, 
    17316, 
    17319, 
    17322, 
    17325, 
    17328, 
    17331, 
    17334, 
    17337, 
    17340, 
    17343, 
    17346, 
    17349, 
    17352, 
    17355, 
    17358, 
    17361, 
    17364, 
    17367, 
    17370, 
    17373, 
    17376, 
    17379, 
    17382, 
    17385, 
    17388, 
    17391, 
    17394, 
    17397, 
    17400, 
    17403, 
    17406, 
    17409, 
    17412, 
    17415, 
    17418, 
    17421, 
    17424, 
    17427, 
    17430, 
    17433, 
    17436, 
    17439, 
    17442, 
    17445, 
    17448, 
    17451, 
    17454, 
    17457, 
    17460, 
    17463, 
    17466, 
    17469, 
    17472, 
    17475, 
    17478, 
    17481, 
    17484, 
    17487, 
    17490, 
    17493, 
    17496, 
    17499, 
    17502, 
    17505, 
    17508, 
    17511, 
    17514, 
    17517, 
    17520, 
    17523, 
    17526, 
    17529, 
    17532, 
    17535, 
    17538, 
    17541, 
    17544, 
    17547, 
    17550, 
    17553, 
    17556, 
    17559, 
    17562, 
    17565, 
    17568, 
    17571, 
    17574, 
    17577, 
    17580, 
    17583, 
    17586, 
    17589, 
    17592, 
    17595, 
    17598, 
    17601, 
    17604, 
    17607, 
    17610, 
    17613, 
    17616, 
    17619, 
    17622, 
    17625, 
    17628, 
    17631, 
    17634, 
    17637, 
    17640, 
    17643, 
    17646, 
    17649, 
    17652, 
    17655, 
    17658, 
    17661, 
    17664, 
    17667, 
    17670, 
    17673, 
    17676, 
    17679, 
    17682, 
    17685, 
    17688, 
    17691, 
    17694, 
    17697, 
    17700, 
    17703, 
    17706, 
    17709, 
    17712, 
    17715, 
    17718, 
    17721, 
    17724, 
    17727, 
    17730, 
    17733, 
    17736, 
    17739, 
    17742, 
    17745, 
    17748, 
    17751, 
    17754, 
    17757, 
    17760, 
    17763, 
    17766, 
    17769, 
    17772, 
    17775, 
    17778, 
    17781, 
    17784, 
    17787, 
    17790, 
    17793, 
    17796, 
    17799, 
    17802, 
    17805, 
    17808, 
    17811, 
    17814, 
    17817, 
    17820, 
    17823, 
    17826, 
    17829, 
    17832, 
    17835, 
    17838, 
    17841, 
    17844, 
    17847, 
    17850, 
    17853, 
    17856, 
    17859, 
    17862, 
    17865, 
    17868, 
    17871, 
    17874, 
    17877, 
    17880, 
    17883, 
    17886, 
    17889, 
    17892, 
    17895, 
    17898, 
    17901, 
    17904, 
    17907, 
    17910, 
    17913, 
    17916, 
    17919, 
    17922, 
    17925, 
    17928, 
    17931, 
    17934, 
    17937, 
    17940, 
    17943, 
    17946, 
    17949, 
    17952, 
    17955, 
    17958, 
    17961, 
    17964, 
    17967, 
    17970, 
    17973, 
    17976, 
    17979, 
    17982, 
    17985, 
    17988, 
    17991, 
    17994, 
    17997, 
    18000, 
    18003, 
    18006, 
    18009, 
    18012, 
    18015, 
    18018, 
    18021, 
    18024, 
    18027, 
    18030, 
    18033, 
    18036, 
    18039, 
    18042, 
    18045, 
    18048, 
    18051, 
    18054, 
    18057, 
    18060, 
    18063, 
    18066, 
    18069, 
    18072, 
    18075, 
    18078, 
    18081, 
    18084, 
    18087, 
    18090, 
    18093, 
    18096, 
    18099, 
    18102, 
    18105, 
    18108, 
    18111, 
    18114, 
    18117, 
    18120, 
    18123, 
    18126, 
    18129, 
    18132, 
    18135, 
    18138, 
    18141, 
    18144, 
    18147, 
    18150, 
    18153, 
    18156, 
    18159, 
    18162, 
    18165, 
    18168, 
    18171, 
    18174, 
    18177, 
    18180, 
    18183, 
    18186, 
    18189, 
    18192, 
    18195, 
    18198, 
    18201, 
    18204, 
    18207, 
    18210, 
    18213, 
    18216, 
    18219, 
    18222, 
    18225, 
    18228, 
    18231, 
    18234, 
    18237, 
    18240, 
    18243, 
    18246, 
    18249, 
    18252, 
    18255, 
    18258, 
    18261, 
    18264, 
    18267, 
    18270, 
    18273, 
    18276, 
    18279, 
    18282, 
    18285, 
    18288, 
    18291, 
    18294, 
    18297, 
    18300, 
    18303, 
    18306, 
    18309, 
    18312, 
    18315, 
    18318, 
    18321, 
    18324, 
    18327, 
    18330, 
    18333, 
    18336, 
    18339, 
    18342, 
    18345, 
    18348, 
    18351, 
    18354, 
    18357, 
    18360, 
    18363, 
    18366, 
    18369, 
    18372, 
    18375, 
    18378, 
    18381, 
    18384, 
    18387, 
    18390, 
    18393, 
    18396, 
    18399, 
    18402, 
    18405, 
    18408, 
    18411, 
    18414, 
    18417, 
    18420, 
    18423, 
    18426, 
    18429, 
    18432, 
    18435, 
    18438, 
    18441, 
    18444, 
    18447, 
    18450, 
    18453, 
    18456, 
    18459, 
    18462, 
    18465, 
    18468, 
    18471, 
    18474, 
    18477, 
    18480, 
    18483, 
    18486, 
    18489, 
    18492, 
    18495, 
    18498, 
    18501, 
    18504, 
    18507, 
    18510, 
    18513, 
    18516, 
    18519, 
    18522, 
    18525, 
    18528, 
    18531, 
    18534, 
    18537, 
    18540, 
    18543, 
    18546, 
    18549, 
    18552, 
    18555, 
    18558, 
    18561, 
    18564, 
    18567, 
    18570, 
    18573, 
    18576, 
    18579, 
    18582, 
    18585, 
    18588, 
    18591, 
    18594, 
    18597, 
    18600, 
    18603, 
    18606, 
    18609, 
    18612, 
    18615, 
    18618, 
    18621, 
    18624, 
    18627, 
    18630, 
    18633, 
    18636, 
    18639, 
    18642, 
    18645, 
    18648, 
    18651, 
    18654, 
    18657, 
    18660, 
    18663, 
    18666, 
    18669, 
    18672, 
    18675, 
    18678, 
    18681, 
    18684, 
    18687, 
    18690, 
    18693, 
    18696, 
    18699, 
    18702, 
    18705, 
    18708, 
    18711, 
    18714, 
    18717, 
    18720, 
    18723, 
    18726, 
    18729, 
    18732, 
    18735, 
    18738, 
    18741, 
    18744, 
    18747, 
    18750, 
    18753, 
    18756, 
    18759, 
    18762, 
    18765, 
    18768, 
    18771, 
    18774, 
    18777, 
    18780, 
    18783, 
    18786, 
    18789, 
    18792, 
    18795, 
    18798, 
    18801, 
    18804, 
    18807, 
    18810, 
    18813, 
    18816, 
    18819, 
    18822, 
    18825, 
    18828, 
    18831, 
    18834, 
    18837, 
    18840, 
    18843, 
    18846, 
    18849, 
    18852, 
    18855, 
    18858, 
    18861, 
    18864, 
    18867, 
    18870, 
    18873, 
    18876, 
    18879, 
    18882, 
    18885, 
    18888, 
    18891, 
    18894, 
    18897, 
    18900, 
    18903, 
    18906, 
    18909, 
    18912, 
    18915, 
    18918, 
    18921, 
    18924, 
    18927, 
    18930, 
    18933, 
    18936, 
    18939, 
    18942, 
    18945, 
    18948, 
    18951, 
    18954, 
    18957, 
    18960, 
    18963, 
    18966, 
    18969, 
    18972, 
    18975, 
    18978, 
    18981, 
    18984, 
    18987, 
    18990, 
    18993, 
    18996, 
    18999, 
    19002, 
    19005, 
    19008, 
    19011, 
    19014, 
    19017, 
    19020, 
    19023, 
    19026, 
    19029, 
    19032, 
    19035, 
    19038, 
    19041, 
    19044, 
    19047, 
    19050, 
    19053, 
    19056, 
    19059, 
    19062, 
    19065, 
    19068, 
    19071, 
    19074, 
    19077, 
    19080, 
    19083, 
    19086, 
    19089, 
    19092, 
    19095, 
    19098, 
    19101, 
    19104, 
    19107, 
    19110, 
    19113, 
    19116, 
    19119, 
    19122, 
    19125, 
    19128, 
    19131, 
    19134, 
    19137, 
    19140, 
    19143, 
    19146, 
    19149, 
    19152, 
    19155, 
    19158, 
    19161, 
    19164, 
    19167, 
    19170, 
    19173, 
    19176, 
    19179, 
    19182, 
    19185, 
    19188, 
    19191, 
    19194, 
    19197, 
    19200, 
    19203, 
    19206, 
    19209, 
    19212, 
    19215, 
    19218, 
    19221, 
    19224, 
    19227, 
    19230, 
    19233, 
    19236, 
    19239, 
    19242, 
    19245, 
    19248, 
    19251, 
    19254, 
    19257, 
    19260, 
    19263, 
    19266, 
    19269, 
    19272, 
    19275, 
    19278, 
    19281, 
    19284, 
    19287, 
    19290, 
    19293, 
    19296, 
    19299, 
    19302, 
    19305, 
    19308, 
    19311, 
    19314, 
    19317, 
    19320, 
    19323, 
    19326, 
    19329, 
    19332, 
    19335, 
    19338, 
    19341, 
    19344, 
    19347, 
    19350, 
    19353, 
    19356, 
    19359, 
    19362, 
    19365, 
    19368, 
    19371, 
    19374, 
    19377, 
    19380, 
    19383, 
    19386, 
    19389, 
    19392, 
    19395, 
    19398, 
    19401, 
    19404, 
    19407, 
    19410, 
    19413, 
    19416, 
    19419, 
    19422, 
    19425, 
    19428, 
    19431, 
    19434, 
    19437, 
    19440, 
    19443, 
    19446, 
    19449, 
    19452, 
    19455, 
    19458, 
    19461, 
    19464, 
    19467, 
    19470, 
    19473, 
    19476, 
    19479, 
    19482, 
    19485, 
    19488, 
    19491, 
    19494, 
    19497, 
    19500, 
    19503, 
    19506, 
    19509, 
    19512, 
    19515, 
    19518, 
    19521, 
    19524, 
    19527, 
    19530, 
    19533, 
    19536, 
    19539, 
    19542, 
    19545, 
    19548, 
    19551, 
    19554, 
    19557, 
    19560, 
    19563, 
    19566, 
    19569, 
    19572, 
    19575, 
    19578, 
    19581, 
    19584, 
    19587, 
    19590, 
    19593, 
    19596, 
    19599, 
    19602, 
    19605, 
    19608, 
    19611, 
    19614, 
    19617, 
    19620, 
    19623, 
    19626, 
    19629, 
    19632, 
    19635, 
    19638, 
    19641, 
    19644, 
    19647, 
    19650, 
    19653, 
    19656, 
    19659, 
    19662, 
    19665, 
    19668, 
    19671, 
    19674, 
    19677, 
    19680, 
    19683, 
    19686, 
    19689, 
    19692, 
    19695, 
    19698, 
    19701, 
    19704, 
    19707, 
    19710, 
    19713, 
    19716, 
    19719, 
    19722, 
    19725, 
    19728, 
    19731, 
    19734, 
    19737, 
    19740, 
    19743, 
    19746, 
    19749, 
    19752, 
    19755, 
    19758, 
    19761, 
    19764, 
    19767, 
    19770, 
    19773, 
    19776, 
    19779, 
    19782, 
    19785, 
    19788, 
    19791, 
    19794, 
    19797, 
    19800, 
    19803, 
    19806, 
    19809, 
    19812, 
    19815, 
    19818, 
    19821, 
    19824, 
    19827, 
    19830, 
    19833, 
    19836, 
    19839, 
    19842, 
    19845, 
    19848, 
    19851, 
    19854, 
    19857, 
    19860, 
    19863, 
    19866, 
    19869, 
    19872, 
    19875, 
    19878, 
    19881, 
    19884, 
    19887, 
    19890, 
    19893, 
    19896, 
    19899, 
    19902, 
    19905, 
    19908, 
    19911, 
    19914, 
    19917, 
    19920, 
    19923, 
    19926, 
    19929, 
    19932, 
    19935, 
    19938, 
    19941, 
    19944, 
    19947, 
    19950, 
    19953, 
    19956, 
    19959, 
    19962, 
    19965, 
    19968, 
    19971, 
    19974, 
    19977, 
    19980, 
    19983, 
    19986, 
    19989, 
    19992, 
    19995, 
    19998, 
    20001, 
    20004, 
    20007, 
    20010, 
    20013, 
    20016, 
    20019, 
    20022, 
    20025, 
    20028, 
    20031, 
    20034, 
    20037, 
    20040, 
    20043, 
    20046, 
    20049, 
    20052, 
    20055, 
    20058, 
    20061, 
    20064, 
    20067, 
    20070, 
    20073, 
    20076, 
    20079, 
    20082, 
    20085, 
    20088, 
    20091, 
    20094, 
    20097, 
    20100, 
    20103, 
    20106, 
    20109, 
    20112, 
    20115, 
    20118, 
    20121, 
    20124, 
    20127, 
    20130, 
    20133, 
    20136, 
    20139, 
    20142, 
    20145, 
    20148, 
    20151, 
    20154, 
    20157, 
    20160, 
    20163, 
    20166, 
    20169, 
    20172, 
    20175, 
    20178, 
    20181, 
    20184, 
    20187, 
    20190, 
    20193, 
    20196, 
    20199, 
    20202, 
    20205, 
    20208, 
    20211, 
    20214, 
    20217, 
    20220, 
    20223, 
    20226, 
    20229, 
    20232, 
    20235, 
    20238, 
    20241, 
    20244, 
    20247, 
    20250, 
    20253, 
    20256, 
    20259, 
    20262, 
    20265, 
    20268, 
    20271, 
    20274, 
    20277, 
    20280, 
    20283, 
    20286, 
    20289, 
    20292, 
    20295, 
    20298, 
    20301, 
    20304, 
    20307, 
    20310, 
    20313, 
    20316, 
    20319, 
    20322, 
    20325, 
    20328, 
    20331, 
    20334, 
    20337, 
    20340, 
    20343, 
    20346, 
    20349, 
    20352, 
    20355, 
    20358, 
    20361, 
    20364, 
    20367, 
    20370, 
    20373, 
    20376, 
    20379, 
    20382, 
    20385, 
    20388, 
    20391, 
    20394, 
    20397, 
    20400, 
    20403, 
    20406, 
    20409, 
    20412, 
    20415, 
    20418, 
    20421, 
    20424, 
    20427, 
    20430, 
    20433, 
    20436, 
    20439, 
    20442, 
    20445, 
    20448, 
    20451, 
    20454, 
    20457, 
    20460, 
    20463, 
    20466, 
    20469, 
    20472, 
    20475, 
    20478, 
    20481, 
    20484, 
    20487, 
    20490, 
    20493, 
    20496, 
    20499, 
    20502, 
    20505, 
    20508, 
    20511, 
    20514, 
    20517, 
    20520, 
    20523, 
    20526, 
    20529, 
    20532, 
    20535, 
    20538, 
    20541, 
    20544, 
    20547, 
    20550, 
    20553, 
    20556, 
    20559, 
    20562, 
    20565, 
    20568, 
    20571, 
    20574, 
    20577, 
    20580, 
    20583, 
    20586, 
    20589, 
    20592, 
    20595, 
    20598, 
    20601, 
    20604, 
    20607, 
    20610, 
    20613, 
    20616, 
    20619, 
    20622, 
    20625, 
    20628, 
    20631, 
    20634, 
    20637, 
    20640, 
    20643, 
    20646, 
    20649, 
    20652, 
    20655, 
    20658, 
    20661, 
    20664, 
    20667, 
    20670, 
    20673, 
    20676, 
    20679, 
    20682, 
    20685, 
    20688, 
    20691, 
    20694, 
    20697, 
    20700, 
    20703, 
    20706, 
    20709, 
    20712, 
    20715, 
    20718, 
    20721, 
    20724, 
    20727, 
    20730, 
    20733, 
    20736, 
    20739, 
    20742, 
    20745, 
    20748, 
    20751, 
    20754, 
    20757, 
    20760, 
    20763, 
    20766, 
    20769, 
    20772, 
    20775, 
    20778, 
    20781, 
    20784, 
    20787, 
    20790, 
    20793, 
    20796, 
    20799, 
    20802, 
    20805, 
    20808, 
    20811, 
    20814, 
    20817, 
    20820, 
    20823, 
    20826, 
    20829, 
    20832, 
    20835, 
    20838, 
    20841, 
    20844, 
    20847, 
    20850, 
    20853, 
    20856, 
    20859, 
    20862, 
    20865, 
    20868, 
    20871, 
    20874, 
    20877, 
    20880, 
    20883, 
    20886, 
    20889, 
    20892, 
    20895, 
    20898, 
    20901, 
    20904, 
    20907, 
    20910, 
    20913, 
    20916, 
    20919, 
    20922, 
    20925, 
    20928, 
    20931, 
    20934, 
    20937, 
    20940, 
    20943, 
    20946, 
    20949, 
    20952, 
    20955, 
    20958, 
    20961, 
    20964, 
    20967, 
    20970, 
    20973, 
    20976, 
    20979, 
    20982, 
    20985, 
    20988, 
    20991, 
    20994, 
    20997, 
    21000, 
    21003, 
    21006, 
    21009, 
    21012, 
    21015, 
    21018, 
    21021, 
    21024, 
    21027, 
    21030, 
    21033, 
    21036, 
    21039, 
    21042, 
    21045, 
    21048, 
    21051, 
    21054, 
    21057, 
    21060, 
    21063, 
    21066, 
    21069, 
    21072, 
    21075, 
    21078, 
    21081, 
    21084, 
    21087, 
    21090, 
    21093, 
    21096, 
    21099, 
    21102, 
    21105, 
    21108, 
    21111, 
    21114, 
    21117, 
    21120, 
    21123, 
    21126, 
    21129, 
    21132, 
    21135, 
    21138, 
    21141, 
    21144, 
    21147, 
    21150, 
    21153, 
    21156, 
    21159, 
    21162, 
    21165, 
    21168, 
    21171, 
    21174, 
    21177, 
    21180, 
    21183, 
    21186, 
    21189, 
    21192, 
    21195, 
    21198, 
    21201, 
    21204, 
    21207, 
    21210, 
    21213, 
    21216, 
    21219, 
    21222, 
    21225, 
    21228, 
    21231, 
    21234, 
    21237, 
    21240, 
    21243, 
    21246, 
    21249, 
    21252, 
    21255, 
    21258, 
    21261, 
    21264, 
    21267, 
    21270, 
    21273, 
    21276, 
    21279, 
    21282, 
    21285, 
    21288, 
    21291, 
    21294, 
    21297, 
    21300, 
    21303, 
    21306, 
    21309, 
    21312, 
    21315, 
    21318, 
    21321, 
    21324, 
    21327, 
    21330, 
    21333, 
    21336, 
    21339, 
    21342, 
    21345, 
    21348, 
    21351, 
    21354, 
    21357, 
    21360, 
    21363, 
    21366, 
    21369, 
    21372, 
    21375, 
    21378, 
    21381, 
    21384, 
    21387, 
    21390, 
    21393, 
    21396, 
    21399, 
    21402, 
    21405, 
    21408, 
    21411, 
    21414, 
    21417, 
    21420, 
    21423, 
    21426, 
    21429, 
    21432, 
    21435, 
    21438, 
    21441, 
    21444, 
    21447, 
    21450, 
    21453, 
    21456, 
    21459, 
    21462, 
    21465, 
    21468, 
    21471, 
    21474, 
    21477, 
    21480, 
    21483, 
    21486, 
    21489, 
    21492, 
    21495, 
    21498, 
    21501, 
    21504, 
    21507, 
    21510, 
    21513, 
    21516, 
    21519, 
    21522, 
    21525, 
    21528, 
    21531, 
    21534, 
    21537, 
    21540, 
    21543, 
    21546, 
    21549, 
    21552, 
    21555, 
    21558, 
    21561, 
    21564, 
    21567, 
    21570, 
    21573, 
    21576, 
    21579, 
    21582, 
    21585, 
    21588, 
    21591, 
    21594, 
    21597, 
    21600, 
    21603, 
    21606, 
    21609, 
    21612, 
    21615, 
    21618, 
    21621, 
    21624, 
    21627, 
    21630, 
    21633, 
    21636, 
    21639, 
    21642, 
    21645, 
    21648, 
    21651, 
    21654, 
    21657, 
    21660, 
    21663, 
    21666, 
    21669, 
    21672, 
    21675, 
    21678, 
    21681, 
    21684, 
    21687, 
    21690, 
    21693, 
    21696, 
    21699, 
    21702, 
    21705, 
    21708, 
    21711, 
    21714, 
    21717, 
    21720, 
    21723, 
    21726, 
    21729, 
    21732, 
    21735, 
    21738, 
    21741, 
    21744, 
    21747, 
    21750, 
    21753, 
    21756, 
    21759, 
    21762, 
    21765, 
    21768, 
    21771, 
    21774, 
    21777, 
    21780, 
    21783, 
    21786, 
    21789, 
    21792, 
    21795, 
    21798, 
    21801, 
    21804, 
    21807, 
    21810, 
    21813, 
    21816, 
    21819, 
    21822, 
    21825, 
    21828, 
    21831, 
    21834, 
    21837, 
    21840, 
    21843, 
    21846, 
    21849, 
    21852, 
    21855, 
    21858, 
    21861, 
    21864, 
    21867, 
    21870, 
    21873, 
    21876, 
    21879, 
    21882, 
    21885, 
    21888, 
    21891, 
    21894, 
    21897, 
    21900, 
    21903, 
    21906, 
    21909, 
    21912, 
    21915, 
    21918, 
    21921, 
    21924, 
    21927, 
    21930, 
    21933, 
    21936, 
    21939, 
    21942, 
    21945, 
    21948, 
    21951, 
    21954, 
    21957, 
    21960, 
    21963, 
    21966, 
    21969, 
    21972, 
    21975, 
    21978, 
    21981, 
    21984, 
    21987, 
    21990, 
    21993, 
    21996, 
    21999, 
    22002, 
    22005, 
    22008, 
    22011, 
    22014, 
    22017, 
    22020, 
    22023, 
    22026, 
    22029, 
    22032, 
    22035, 
    22038, 
    22041, 
    22044, 
    22047, 
    22050, 
    22053, 
    22056, 
    22059, 
    22062, 
    22065, 
    22068, 
    22071, 
    22074, 
    22077, 
    22080, 
    22083, 
    22086, 
    22089, 
    22092, 
    22095, 
    22098, 
    22101, 
    22104, 
    22107, 
    22110, 
    22113, 
    22116, 
    22119, 
    22122, 
    22125, 
    22128, 
    22131, 
    22134, 
    22137, 
    22140, 
    22143, 
    22146, 
    22149, 
    22152, 
    22155, 
    22158, 
    22161, 
    22164, 
    22167, 
    22170, 
    22173, 
    22176, 
    22179, 
    22182, 
    22185, 
    22188, 
    22191, 
    22194, 
    22197, 
    22200, 
    22203, 
    22206, 
    22209, 
    22212, 
    22215, 
    22218, 
    22221, 
    22224, 
    22227, 
    22230, 
    22233, 
    22236, 
    22239, 
    22242, 
    22245, 
    22248, 
    22251, 
    22254, 
    22257, 
    22260, 
    22263, 
    22266, 
    22269, 
    22272, 
    22275, 
    22278, 
    22281, 
    22284, 
    22287, 
    22290, 
    22293, 
    22296, 
    22299, 
    22302, 
    22305, 
    22308, 
    22311, 
    22314, 
    22317, 
    22320, 
    22323, 
    22326, 
    22329, 
    22332, 
    22335, 
    22338, 
    22341, 
    22344, 
    22347, 
    22350, 
    22353, 
    22356, 
    22359, 
    22362, 
    22365, 
    22368, 
    22371, 
    22374, 
    22377, 
    22380, 
    22383, 
    22386, 
    22389, 
    22392, 
    22395, 
    22398, 
    22401, 
    22404, 
    22407, 
    22410, 
    22413, 
    22416, 
    22419, 
    22422, 
    22425, 
    22428, 
    22431, 
    22434, 
    22437, 
    22440, 
    22443, 
    22446, 
    22449, 
    22452, 
    22455, 
    22458, 
    22461, 
    22464, 
    22467, 
    22470, 
    22473, 
    22476, 
    22479, 
    22482, 
    22485, 
    22488, 
    22491, 
    22494, 
    22497, 
    22500, 
    22503, 
    22506, 
    22509, 
    22512, 
    22515, 
    22518, 
    22521, 
    22524, 
    22527, 
    22530, 
    22533, 
    22536, 
    22539, 
    22542, 
    22545, 
    22548, 
    22551, 
    22554, 
    22557, 
    22560, 
    22563, 
    22566, 
    22569, 
    22572, 
    22575, 
    22578, 
    22581, 
    22584, 
    22587, 
    22590, 
    22593, 
    22596, 
    22599, 
    22602, 
    22605, 
    22608, 
    22611, 
    22614, 
    22617, 
    22620, 
    22623, 
    22626, 
    22629, 
    22632, 
    22635, 
    22638, 
    22641, 
    22644, 
    22647, 
    22650, 
    22653, 
    22656, 
    22659, 
    22662, 
    22665, 
    22668, 
    22671, 
    22674, 
    22677, 
    22680, 
    22683, 
    22686, 
    22689, 
    22692, 
    22695, 
    22698, 
    22701, 
    22704, 
    22707, 
    22710, 
    22713, 
    22716, 
    22719, 
    22722, 
    22725, 
    22728, 
    22731, 
    22734, 
    22737, 
    22740, 
    22743, 
    22746, 
    22749, 
    22752, 
    22755, 
    22758, 
    22761, 
    22764, 
    22767, 
    22770, 
    22773, 
    22776, 
    22779, 
    22782, 
    22785, 
    22788, 
    22791, 
    22794, 
    22797, 
    22800, 
    22803, 
    22806, 
    22809, 
    22812, 
    22815, 
    22818, 
    22821, 
    22824, 
    22827, 
    22830, 
    22833, 
    22836, 
    22839, 
    22842, 
    22845, 
    22848, 
    22851, 
    22854, 
    22857, 
    22860, 
    22863, 
    22866, 
    22869, 
    22872, 
    22875, 
    22878, 
    22881, 
    22884, 
    22887, 
    22890, 
    22893, 
    22896, 
    22899, 
    22902, 
    22905, 
    22908, 
    22911, 
    22914, 
    22917, 
    22920, 
    22923, 
    22926, 
    22929, 
    22932, 
    22935, 
    22938, 
    22941, 
    22944, 
    22947, 
    22950, 
    22953, 
    22956, 
    22959, 
    22962, 
    22965, 
    22968, 
    22971, 
    22974, 
    22977, 
    22980, 
    22983, 
    22986, 
    22989, 
    22992, 
    22995, 
    22998, 
    23001, 
    23004, 
    23007, 
    23010, 
    23013, 
    23016, 
    23019, 
    23022, 
    23025, 
    23028, 
    23031, 
    23034, 
    23037, 
    23040, 
    23043, 
    23046, 
    23049, 
    23052, 
    23055, 
    23058, 
    23061, 
    23064, 
    23067, 
    23070, 
    23073, 
    23076, 
    23079, 
    23082, 
    23085, 
    23088, 
    23091, 
    23094, 
    23097, 
    23100, 
    23103, 
    23106, 
    23109, 
    23112, 
    23115, 
    23118, 
    23121, 
    23124, 
    23127, 
    23130, 
    23133, 
    23136, 
    23139, 
    23142, 
    23145, 
    23148, 
    23151, 
    23154, 
    23157, 
    23160, 
    23163, 
    23166, 
    23169, 
    23172, 
    23175, 
    23178, 
    23181, 
    23184, 
    23187, 
    23190, 
    23193, 
    23196, 
    23199, 
    23202, 
    23205, 
    23208, 
    23211, 
    23214, 
    23217, 
    23220, 
    23223, 
    23226, 
    23229, 
    23232, 
    23235, 
    23238, 
    23241, 
    23244, 
    23247, 
    23250, 
    23253, 
    23256, 
    23259, 
    23262, 
    23265, 
    23268, 
    23271, 
    23274, 
    23277, 
    23280, 
    23283, 
    23286, 
    23289, 
    23292, 
    23295, 
    23298, 
    23301, 
    23304, 
    23307, 
    23310, 
    23313, 
    23316, 
    23319, 
    23322, 
    23325, 
    23328, 
    23331, 
    23334, 
    23337, 
    23340, 
    23343, 
    23346, 
    23349, 
    23352, 
    23355, 
    23358, 
    23361, 
    23364, 
    23367, 
    23370, 
    23373, 
    23376, 
    23379, 
    23382, 
    23385, 
    23388, 
    23391, 
    23394, 
    23397, 
    23400, 
    23403, 
    23406, 
    23409, 
    23412, 
    23415, 
    23418, 
    23421, 
    23424, 
    23427, 
    23430, 
    23433, 
    23436, 
    23439, 
    23442, 
    23445, 
    23448, 
    23451, 
    23454, 
    23457, 
    23460, 
    23463, 
    23466, 
    23469, 
    23472, 
    23475, 
    23478, 
    23481, 
    23484, 
    23487, 
    23490, 
    23493, 
    23496, 
    23499, 
    23502, 
    23505, 
    23508, 
    23511, 
    23514, 
    23517, 
    23520, 
    23523, 
    23526, 
    23529, 
    23532, 
    23535, 
    23538, 
    23541, 
    23544, 
    23547, 
    23550, 
    23553, 
    23556, 
    23559, 
    23562, 
    23565, 
    23568, 
    23571, 
    23574, 
    23577, 
    23580, 
    23583, 
    23586, 
    23589, 
    23592, 
    23595, 
    23598, 
    23601, 
    23604, 
    23607, 
    23610, 
    23613, 
    23616, 
    23619, 
    23622, 
    23625, 
    23628, 
    23631, 
    23634, 
    23637, 
    23640, 
    23643, 
    23646, 
    23649, 
    23652, 
    23655, 
    23658, 
    23661, 
    23664, 
    23667, 
    23670, 
    23673, 
    23676, 
    23679, 
    23682, 
    23685, 
    23688, 
    23691, 
    23694, 
    23697, 
    23700, 
    23703, 
    23706, 
    23709, 
    23712, 
    23715, 
    23718, 
    23721, 
    23724, 
    23727, 
    23730, 
    23733, 
    23736, 
    23739, 
    23742, 
    23745, 
    23748, 
    23751, 
    23754, 
    23757, 
    23760, 
    23763, 
    23766, 
    23769, 
    23772, 
    23775, 
    23778, 
    23781, 
    23784, 
    23787, 
    23790, 
    23793, 
    23796, 
    23799, 
    23802, 
    23805, 
    23808, 
    23811, 
    23814, 
    23817, 
    23820, 
    23823, 
    23826, 
    23829, 
    23832, 
    23835, 
    23838, 
    23841, 
    23844, 
    23847, 
    23850, 
    23853, 
    23856, 
    23859, 
    23862, 
    23865, 
    23868, 
    23871, 
    23874, 
    23877, 
    23880, 
    23883, 
    23886, 
    23889, 
    23892, 
    23895, 
    23898, 
    23901, 
    23904, 
    23907, 
    23910, 
    23913, 
    23916, 
    23919, 
    23922, 
    23925, 
    23928, 
    23931, 
    23934, 
    23937, 
    23940, 
    23943, 
    23946, 
    23949, 
    23952, 
    23955, 
    23958, 
    23961, 
    23964, 
    23967, 
    23970, 
    23973, 
    23976, 
    23979, 
    23982, 
    23985, 
    23988, 
    23991, 
    23994, 
    23997, 
    24000, 
    24003, 
    24006, 
    24009, 
    24012, 
    24015, 
    24018, 
    24021, 
    24024, 
    24027, 
    24030, 
    24033, 
    24036, 
    24039, 
    24042, 
    24045, 
    24048, 
    24051, 
    24054, 
    24057, 
    24060, 
    24063, 
    24066, 
    24069, 
    24072, 
    24075, 
    24078, 
    24081, 
    24084, 
    24087, 
    24090, 
    24093, 
    24096, 
    24099, 
    24102, 
    24105, 
    24108, 
    24111, 
    24114, 
    24117, 
    24120, 
    24123, 
    24126, 
    24129, 
    24132, 
    24135, 
    24138, 
    24141, 
    24144, 
    24147, 
    24150, 
    24153, 
    24156, 
    24159, 
    24162, 
    24165, 
    24168, 
    24171, 
    24174, 
    24177, 
    24180, 
    24183, 
    24186, 
    24189, 
    24192, 
    24195, 
    24198, 
    24201, 
    24204, 
    24207, 
    24210, 
    24213, 
    24216, 
    24219, 
    24222, 
    24225, 
    24228, 
    24231, 
    24234, 
    24237, 
    24240, 
    24243, 
    24246, 
    24249, 
    24252, 
    24255, 
    24258, 
    24261, 
    24264, 
    24267, 
    24270, 
    24273, 
    24276, 
    24279, 
    24282, 
    24285, 
    24288, 
    24291, 
    24294, 
    24297, 
    24300, 
    24303, 
    24306, 
    24309, 
    24312, 
    24315, 
    24318, 
    24321, 
    24324, 
    24327, 
    24330, 
    24333, 
    24336, 
    24339, 
    24342, 
    24345, 
    24348, 
    24351, 
    24354, 
    24357, 
    24360, 
    24363, 
    24366, 
    24369, 
    24372, 
    24375, 
    24378, 
    24381, 
    24384, 
    24387, 
    24390, 
    24393, 
    24396, 
    24399, 
    24402, 
    24405, 
    24408, 
    24411, 
    24414, 
    24417, 
    24420, 
    24423, 
    24426, 
    24429, 
    24432, 
    24435, 
    24438, 
    24441, 
    24444, 
    24447, 
    24450, 
    24453, 
    24456, 
    24459, 
    24462, 
    24465, 
    24468, 
    24471, 
    24474, 
    24477, 
    24480, 
    24483, 
    24486, 
    24489, 
    24492, 
    24495, 
    24498, 
    24501, 
    24504, 
    24507, 
    24510, 
    24513, 
    24516, 
    24519, 
    24522, 
    24525, 
    24528, 
    24531, 
    24534, 
    24537, 
    24540, 
    24543, 
    24546, 
    24549, 
    24552, 
    24555, 
    24558, 
    24561, 
    24564, 
    24567, 
    24570, 
    24573, 
    24576, 
    24579, 
    24582, 
    24585, 
    24588, 
    24591, 
    24594, 
    24597, 
    24600, 
    24603, 
    24606, 
    24609, 
    24612, 
    24615, 
    24618, 
    24621, 
    24624, 
    24627, 
    24630, 
    24633, 
    24636, 
    24639, 
    24642, 
    24645, 
    24648, 
    24651, 
    24654, 
    24657, 
    24660, 
    24663, 
    24666, 
    24669, 
    24672, 
    24675, 
    24678, 
    24681, 
    24684, 
    24687, 
    24690, 
    24693, 
    24696, 
    24699, 
    24702, 
    24705, 
    24708, 
    24711, 
    24714, 
    24717, 
    24720, 
    24723, 
    24726, 
    24729, 
    24732, 
    24735, 
    24738, 
    24741, 
    24744, 
    24747, 
    24750, 
    24753, 
    24756, 
    24759, 
    24762, 
    24765, 
    24768, 
    24771, 
    24774, 
    24777, 
    24780, 
    24783, 
    24786, 
    24789, 
    24792, 
    24795, 
    24798, 
    24801, 
    24804, 
    24807, 
    24810, 
    24813, 
    24816, 
    24819, 
    24822, 
    24825, 
    24828, 
    24831, 
    24834, 
    24837, 
    24840, 
    24843, 
    24846, 
    24849, 
    24852, 
    24855, 
    24858, 
    24861, 
    24864, 
    24867, 
    24870, 
    24873, 
    24876, 
    24879, 
    24882, 
    24885, 
    24888, 
    24891, 
    24894, 
    24897, 
    24900, 
    24903, 
    24906, 
    24909, 
    24912, 
    24915, 
    24918, 
    24921, 
    24924, 
    24927, 
    24930, 
    24933, 
    24936, 
    24939, 
    24942, 
    24945, 
    24948, 
    24951, 
    24954, 
    24957, 
    24960, 
    24963, 
    24966, 
    24969, 
    24972, 
    24975, 
    24978, 
    24981, 
    24984, 
    24987, 
    24990, 
    24993, 
    24996, 
    24999, 
    25002, 
    25005, 
    25008, 
    25011, 
    25014, 
    25017, 
    25020, 
    25023, 
    25026, 
    25029, 
    25032, 
    25035, 
    25038, 
    25041, 
    25044, 
    25047, 
    25050, 
    25053, 
    25056, 
    25059, 
    25062, 
    25065, 
    25068, 
    25071, 
    25074, 
    25077, 
    25080, 
    25083, 
    25086, 
    25089, 
    25092, 
    25095, 
    25098, 
    25101, 
    25104, 
    25107, 
    25110, 
    25113, 
    25116, 
    25119, 
    25122, 
    25125, 
    25128, 
    25131, 
    25134, 
    25137, 
    25140, 
    25143, 
    25146, 
    25149, 
    25152, 
    25155, 
    25158, 
    25161, 
    25164, 
    25167, 
    25170, 
    25173, 
    25176, 
    25179, 
    25182, 
    25185, 
    25188, 
    25191, 
    25194, 
    25197, 
    25200, 
    25203, 
    25206, 
    25209, 
    25212, 
    25215, 
    25218, 
    25221, 
    25224, 
    25227, 
    25230, 
    25233, 
    25236, 
    25239, 
    25242, 
    25245, 
    25248, 
    25251, 
    25254, 
    25257, 
    25260, 
    25263, 
    25266, 
    25269, 
    25272, 
    25275, 
    25278, 
    25281, 
    25284, 
    25287, 
    25290, 
    25293, 
    25296, 
    25299, 
    25302, 
    25305, 
    25308, 
    25311, 
    25314, 
    25317, 
    25320, 
    25323, 
    25326, 
    25329, 
    25332, 
    25335, 
    25338, 
    25341, 
    25344, 
    25347, 
    25350, 
    25353, 
    25356, 
    25359, 
    25362, 
    25365, 
    25368, 
    25371, 
    25374, 
    25377, 
    25380, 
    25383, 
    25386, 
    25389, 
    25392, 
    25395, 
    25398, 
    25401, 
    25404, 
    25407, 
    25410, 
    25413, 
    25416, 
    25419, 
    25422, 
    25425, 
    25428, 
    25431, 
    25434, 
    25437, 
    25440, 
    25443, 
    25446, 
    25449, 
    25452, 
    25455, 
    25458, 
    25461, 
    25464, 
    25467, 
    25470, 
    25473, 
    25476, 
    25479, 
    25482, 
    25485, 
    25488, 
    25491, 
    25494, 
    25497, 
    25500, 
    25503, 
    25506, 
    25509, 
    25512, 
    25515, 
    25518, 
    25521, 
    25524, 
    25527, 
    25530, 
    25533, 
    25536, 
    25539, 
    25542, 
    25545, 
    25548, 
    25551, 
    25554, 
    25557, 
    25560, 
    25563, 
    25566, 
    25569, 
    25572, 
    25575, 
    25578, 
    25581, 
    25584, 
    25587, 
    25590, 
    25593, 
    25596, 
    25599, 
    25602, 
    25605, 
    25608, 
    25611, 
    25614, 
    25617, 
    25620, 
    25623, 
    25626, 
    25629, 
    25632, 
    25635, 
    25638, 
    25641, 
    25644, 
    25647, 
    25650, 
    25653, 
    25656, 
    25659, 
    25662, 
    25665, 
    25668, 
    25671, 
    25674, 
    25677, 
    25680, 
    25683, 
    25686, 
    25689, 
    25692, 
    25695, 
    25698, 
    25701, 
    25704, 
    25707, 
    25710, 
    25713, 
    25716, 
    25719, 
    25722, 
    25725, 
    25728, 
    25731, 
    25734, 
    25737, 
    25740, 
    25743, 
    25746, 
    25749, 
    25752, 
    25755, 
    25758, 
    25761, 
    25764, 
    25767, 
    25770, 
    25773, 
    25776, 
    25779, 
    25782, 
    25785, 
    25788, 
    25791, 
    25794, 
    25797, 
    25800, 
    25803, 
    25806, 
    25809, 
    25812, 
    25815, 
    25818, 
    25821, 
    25824, 
    25827, 
    25830, 
    25833, 
    25836, 
    25839, 
    25842, 
    25845, 
    25848, 
    25851, 
    25854, 
    25857, 
    25860, 
    25863, 
    25866, 
    25869, 
    25872, 
    25875, 
    25878, 
    25881, 
    25884, 
    25887, 
    25890, 
    25893, 
    25896, 
    25899, 
    25902, 
    25905, 
    25908, 
    25911, 
    25914, 
    25917, 
    25920, 
    25923, 
    25926, 
    25929, 
    25932, 
    25935, 
    25938, 
    25941, 
    25944, 
    25947, 
    25950, 
    25953, 
    25956, 
    25959, 
    25962, 
    25965, 
    25968, 
    25971, 
    25974, 
    25977, 
    25980, 
    25983, 
    25986, 
    25989, 
    25992, 
    25995, 
    25998, 
    26001, 
    26004, 
    26007, 
    26010, 
    26013, 
    26016, 
    26019, 
    26022, 
    26025, 
    26028, 
    26031, 
    26034, 
    26037, 
    26040, 
    26043, 
    26046, 
    26049, 
    26052, 
    26055, 
    26058, 
    26061, 
    26064, 
    26067, 
    26070, 
    26073, 
    26076, 
    26079, 
    26082, 
    26085, 
    26088, 
    26091, 
    26094, 
    26097, 
    26100, 
    26103, 
    26106, 
    26109, 
    26112, 
    26115, 
    26118, 
    26121, 
    26124, 
    26127, 
    26130, 
    26133, 
    26136, 
    26139, 
    26142, 
    26145, 
    26148, 
    26151, 
    26154, 
    26157, 
    26160, 
    26163, 
    26166, 
    26169, 
    26172, 
    26175, 
    26178, 
    26181, 
    26184, 
    26187, 
    26190, 
    26193, 
    26196, 
    26199, 
    26202, 
    26205, 
    26208, 
    26211, 
    26214, 
    26217, 
    26220, 
    26223, 
    26226, 
    26229, 
    26232, 
    26235, 
    26238, 
    26241, 
    26244, 
    26247, 
    26250, 
    26253, 
    26256, 
    26259, 
    26262, 
    26265, 
    26268, 
    26271, 
    26274, 
    26277, 
    26280, 
    26283, 
    26286, 
    26289, 
    26292, 
    26295, 
    26298, 
    26301, 
    26304, 
    26307, 
    26310, 
    26313, 
    26316, 
    26319, 
    26322, 
    26325, 
    26328, 
    26331, 
    26334, 
    26337, 
    26340, 
    26343, 
    26346, 
    26349, 
    26352, 
    26355, 
    26358, 
    26361, 
    26364, 
    26367, 
    26370, 
    26373, 
    26376, 
    26379, 
    26382, 
    26385, 
    26388, 
    26391, 
    26394, 
    26397, 
    26400, 
    26403, 
    26406, 
    26409, 
    26412, 
    26415, 
    26418, 
    26421, 
    26424, 
    26427, 
    26430, 
    26433, 
    26436, 
    26439, 
    26442, 
    26445, 
    26448, 
    26451, 
    26454, 
    26457, 
    26460, 
    26463, 
    26466, 
    26469, 
    26472, 
    26475, 
    26478, 
    26481, 
    26484, 
    26487, 
    26490, 
    26493, 
    26496, 
    26499, 
    26502, 
    26505, 
    26508, 
    26511, 
    26514, 
    26517, 
    26520, 
    26523, 
    26526, 
    26529, 
    26532, 
    26535, 
    26538, 
    26541, 
    26544, 
    26547, 
    26550, 
    26553, 
    26556, 
    26559, 
    26562, 
    26565, 
    26568, 
    26571, 
    26574, 
    26577, 
    26580, 
    26583, 
    26586, 
    26589, 
    26592, 
    26595, 
    26598, 
    26601, 
    26604, 
    26607, 
    26610, 
    26613, 
    26616, 
    26619, 
    26622, 
    26625, 
    26628, 
    26631, 
    26634, 
    26637, 
    26640, 
    26643, 
    26646, 
    26649, 
    26652, 
    26655, 
    26658, 
    26661, 
    26664, 
    26667, 
    26670, 
    26673, 
    26676, 
    26679, 
    26682, 
    26685, 
    26688, 
    26691, 
    26694, 
    26697, 
    26700, 
    26703, 
    26706, 
    26709, 
    26712, 
    26715, 
    26718, 
    26721, 
    26724, 
    26727, 
    26730, 
    26733, 
    26736, 
    26739, 
    26742, 
    26745, 
    26748, 
    26751, 
    26754, 
    26757, 
    26760, 
    26763, 
    26766, 
    26769, 
    26772, 
    26775, 
    26778, 
    26781, 
    26784, 
    26787, 
    26790, 
    26793, 
    26796, 
    26799, 
    26802, 
    26805, 
    26808, 
    26811, 
    26814, 
    26817, 
    26820, 
    26823, 
    26826, 
    26829, 
    26832, 
    26835, 
    26838, 
    26841, 
    26844, 
    26847, 
    26850, 
    26853, 
    26856, 
    26859, 
    26862, 
    26865, 
    26868, 
    26871, 
    26874, 
    26877, 
    26880, 
    26883, 
    26886, 
    26889, 
    26892, 
    26895, 
    26898, 
    26901, 
    26904, 
    26907, 
    26910, 
    26913, 
    26916, 
    26919, 
    26922, 
    26925, 
    26928, 
    26931, 
    26934, 
    26937, 
    26940, 
    26943, 
    26946, 
    26949, 
    26952, 
    26955, 
    26958, 
    26961, 
    26964, 
    26967, 
    26970, 
    26973, 
    26976, 
    26979, 
    26982, 
    26985, 
    26988, 
    26991, 
    26994, 
    26997, 
    27000, 
    27003, 
    27006, 
    27009, 
    27012, 
    27015, 
    27018, 
    27021, 
    27024, 
    27027, 
    27030, 
    27033, 
    27036, 
    27039, 
    27042, 
    27045, 
    27048, 
    27051, 
    27054, 
    27057, 
    27060, 
    27063, 
    27066, 
    27069, 
    27072, 
    27075, 
    27078, 
    27081, 
    27084, 
    27087, 
    27090, 
    27093, 
    27096, 
    27099, 
    27102, 
    27105, 
    27108, 
    27111, 
    27114, 
    27117, 
    27120, 
    27123, 
    27126, 
    27129, 
    27132, 
    27135, 
    27138, 
    27141, 
    27144, 
    27147, 
    27150, 
    27153, 
    27156, 
    27159, 
    27162, 
    27165, 
    27168, 
    27171, 
    27174, 
    27177, 
    27180, 
    27183, 
    27186, 
    27189, 
    27192, 
    27195, 
    27198, 
    27201, 
    27204, 
    27207, 
    27210, 
    27213, 
    27216, 
    27219, 
    27222, 
    27225, 
    27228, 
    27231, 
    27234, 
    27237, 
    27240, 
    27243, 
    27246, 
    27249, 
    27252, 
    27255, 
    27258, 
    27261, 
    27264, 
    27267, 
    27270, 
    27273, 
    27276, 
    27279, 
    27282, 
    27285, 
    27288, 
    27291, 
    27294, 
    27297, 
    27300, 
    27303, 
    27306, 
    27309, 
    27312, 
    27315, 
    27318, 
    27321, 
    27324, 
    27327, 
    27330, 
    27333, 
    27336, 
    27339, 
    27342, 
    27345, 
    27348, 
    27351, 
    27354, 
    27357, 
    27360, 
    27363, 
    27366, 
    27369, 
    27372, 
    27375, 
    27378, 
    27381, 
    27384, 
    27387, 
    27390, 
    27393, 
    27396, 
    27399, 
    27402, 
    27405, 
    27408, 
    27411, 
    27414, 
    27417, 
    27420, 
    27423, 
    27426, 
    27429, 
    27432, 
    27435, 
    27438, 
    27441, 
    27444, 
    27447, 
    27450, 
    27453, 
    27456, 
    27459, 
    27462, 
    27465, 
    27468, 
    27471, 
    27474, 
    27477, 
    27480, 
    27483, 
    27486, 
    27489, 
    27492, 
    27495, 
    27498, 
    27501, 
    27504, 
    27507, 
    27510, 
    27513, 
    27516, 
    27519, 
    27522, 
    27525, 
    27528, 
    27531, 
    27534, 
    27537, 
    27540, 
    27543, 
    27546, 
    27549, 
    27552, 
    27555, 
    27558, 
    27561, 
    27564, 
    27567, 
    27570, 
    27573, 
    27576, 
    27579, 
    27582, 
    27585, 
    27588, 
    27591, 
    27594, 
    27597, 
    27600, 
    27603, 
    27606, 
    27609, 
    27612, 
    27615, 
    27618, 
    27621, 
    27624, 
    27627, 
    27630, 
    27633, 
    27636, 
    27639, 
    27642, 
    27645, 
    27648, 
    27651, 
    27654, 
    27657, 
    27660, 
    27663, 
    27666, 
    27669, 
    27672, 
    27675, 
    27678, 
    27681, 
    27684, 
    27687, 
    27690, 
    27693, 
    27696, 
    27699, 
    27702, 
    27705, 
    27708, 
    27711, 
    27714, 
    27717, 
    27720, 
    27723, 
    27726, 
    27729, 
    27732, 
    27735, 
    27738, 
    27741, 
    27744, 
    27747, 
    27750, 
    27753, 
    27756, 
    27759, 
    27762, 
    27765, 
    27768, 
    27771, 
    27774, 
    27777, 
    27780, 
    27783, 
    27786, 
    27789, 
    27792, 
    27795, 
    27798, 
    27801, 
    27804, 
    27807, 
    27810, 
    27813, 
    27816, 
    27819, 
    27822, 
    27825, 
    27828, 
    27831, 
    27834, 
    27837, 
    27840, 
    27843, 
    27846, 
    27849, 
    27852, 
    27855, 
    27858, 
    27861, 
    27864, 
    27867, 
    27870, 
    27873, 
    27876, 
    27879, 
    27882, 
    27885, 
    27888, 
    27891, 
    27894, 
    27897, 
    27900, 
    27903, 
    27906, 
    27909, 
    27912, 
    27915, 
    27918, 
    27921, 
    27924, 
    27927, 
    27930, 
    27933, 
    27936, 
    27939, 
    27942, 
    27945, 
    27948, 
    27951, 
    27954, 
    27957, 
    27960, 
    27963, 
    27966, 
    27969, 
    27972, 
    27975, 
    27978, 
    27981, 
    27984, 
    27987, 
    27990, 
    27993, 
    27996, 
    27999, 
    28002, 
    28005, 
    28008, 
    28011, 
    28014, 
    28017, 
    28020, 
    28023, 
    28026, 
    28029, 
    28032, 
    28035, 
    28038, 
    28041, 
    28044, 
    28047, 
    28050, 
    28053, 
    28056, 
    28059, 
    28062, 
    28065, 
    28068, 
    28071, 
    28074, 
    28077, 
    28080, 
    28083, 
    28086, 
    28089, 
    28092, 
    28095, 
    28098, 
    28101, 
    28104, 
    28107, 
    28110, 
    28113, 
    28116, 
    28119, 
    28122, 
    28125, 
    28128, 
    28131, 
    28134, 
    28137, 
    28140, 
    28143, 
    28146, 
    28149, 
    28152, 
    28155, 
    28158, 
    28161, 
    28164, 
    28167, 
    28170, 
    28173, 
    28176, 
    28179, 
    28182, 
    28185, 
    28188, 
    28191, 
    28194, 
    28197, 
    28200, 
    28203, 
    28206, 
    28209, 
    28212, 
    28215, 
    28218, 
    28221, 
    28224, 
    28227, 
    28230, 
    28233, 
    28236, 
    28239, 
    28242, 
    28245, 
    28248, 
    28251, 
    28254, 
    28257, 
    28260, 
    28263, 
    28266, 
    28269, 
    28272, 
    28275, 
    28278, 
    28281, 
    28284, 
    28287, 
    28290, 
    28293, 
    28296, 
    28299, 
    28302, 
    28305, 
    28308, 
    28311, 
    28314, 
    28317, 
    28320, 
    28323, 
    28326, 
    28329, 
    28332, 
    28335, 
    28338, 
    28341, 
    28344, 
    28347, 
    28350, 
    28353, 
    28356, 
    28359, 
    28362, 
    28365, 
    28368, 
    28371, 
    28374, 
    28377, 
    28380, 
    28383, 
    28386, 
    28389, 
    28392, 
    28395, 
    28398, 
    28401, 
    28404, 
    28407, 
    28410, 
    28413, 
    28416, 
    28419, 
    28422, 
    28425, 
    28428, 
    28431, 
    28434, 
    28437, 
    28440, 
    28443, 
    28446, 
    28449, 
    28452, 
    28455, 
    28458, 
    28461, 
    28464, 
    28467, 
    28470, 
    28473, 
    28476, 
    28479, 
    28482, 
    28485, 
    28488, 
    28491, 
    28494, 
    28497, 
    28500, 
    28503, 
    28506, 
    28509, 
    28512, 
    28515, 
    28518, 
    28521, 
    28524, 
    28527, 
    28530, 
    28533, 
    28536, 
    28539, 
    28542, 
    28545, 
    28548, 
    28551, 
    28554, 
    28557, 
    28560, 
    28563, 
    28566, 
    28569, 
    28572, 
    28575, 
    28578, 
    28581, 
    28584, 
    28587, 
    28590, 
    28593, 
    28596, 
    28599, 
    28602, 
    28605, 
    28608, 
    28611, 
    28614, 
    28617, 
    28620, 
    28623, 
    28626, 
    28629, 
    28632, 
    28635, 
    28638, 
    28641, 
    28644, 
    28647, 
    28650, 
    28653, 
    28656, 
    28659, 
    28662, 
    28665, 
    28668, 
    28671, 
    28674, 
    28677, 
    28680, 
    28683, 
    28686, 
    28689, 
    28692, 
    28695, 
    28698, 
    28701, 
    28704, 
    28707, 
    28710, 
    28713, 
    28716, 
    28719, 
    28722, 
    28725, 
    28728, 
    28731, 
    28734, 
    28737, 
    28740, 
    28743, 
    28746, 
    28749, 
    28752, 
    28755, 
    28758, 
    28761, 
    28764, 
    28767, 
    28770, 
    28773, 
    28776, 
    28779, 
    28782, 
    28785, 
    28788, 
    28791, 
    28794, 
    28797, 
    28800, 
    28803, 
    28806, 
    28809, 
    28812, 
    28815, 
    28818, 
    28821, 
    28824, 
    28827, 
    28830, 
    28833, 
    28836, 
    28839, 
    28842, 
    28845, 
    28848, 
    28851, 
    28854, 
    28857, 
    28860, 
    28863, 
    28866, 
    28869, 
    28872, 
    28875, 
    28878, 
    28881, 
    28884, 
    28887, 
    28890, 
    28893, 
    28896, 
    28899, 
    28902, 
    28905, 
    28908, 
    28911, 
    28914, 
    28917, 
    28920, 
    28923, 
    28926, 
    28929, 
    28932, 
    28935, 
    28938, 
    28941, 
    28944, 
    28947, 
    28950, 
    28953, 
    28956, 
    28959, 
    28962, 
    28965, 
    28968, 
    28971, 
    28974, 
    28977, 
    28980, 
    28983, 
    28986, 
    28989, 
    28992, 
    28995, 
    28998, 
    29001, 
    29004, 
    29007, 
    29010, 
    29013, 
    29016, 
    29019, 
    29022, 
    29025, 
    29028, 
    29031, 
    29034, 
    29037, 
    29040, 
    29043, 
    29046, 
    29049, 
    29052, 
    29055, 
    29058, 
    29061, 
    29064, 
    29067, 
    29070, 
    29073, 
    29076, 
    29079, 
    29082, 
    29085, 
    29088, 
    29091, 
    29094, 
    29097, 
    29100, 
    29103, 
    29106, 
    29109, 
    29112, 
    29115, 
    29118, 
    29121, 
    29124, 
    29127, 
    29130, 
    29133, 
    29136, 
    29139, 
    29142, 
    29145, 
    29148, 
    29151, 
    29154, 
    29157, 
    29160, 
    29163, 
    29166, 
    29169, 
    29172, 
    29175, 
    29178, 
    29181, 
    29184, 
    29187, 
    29190, 
    29193, 
    29196, 
    29199, 
    29202, 
    29205, 
    29208, 
    29211, 
    29214, 
    29217, 
    29220, 
    29223, 
    29226, 
    29229, 
    29232, 
    29235, 
    29238, 
    29241, 
    29244, 
    29247, 
    29250, 
    29253, 
    29256, 
    29259, 
    29262, 
    29265, 
    29268, 
    29271, 
    29274, 
    29277, 
    29280, 
    29283, 
    29286, 
    29289, 
    29292, 
    29295, 
    29298, 
    29301, 
    29304, 
    29307, 
    29310, 
    29313, 
    29316, 
    29319, 
    29322, 
    29325, 
    29328, 
    29331, 
    29334, 
    29337, 
    29340, 
    29343, 
    29346, 
    29349, 
    29352, 
    29355, 
    29358, 
    29361, 
    29364, 
    29367, 
    29370, 
    29373, 
    29376, 
    29379, 
    29382, 
    29385, 
    29388, 
    29391, 
    29394, 
    29397, 
    29400, 
    29403, 
    29406, 
    29409, 
    29412, 
    29415, 
    29418, 
    29421, 
    29424, 
    29427, 
    29430, 
    29433, 
    29436, 
    29439, 
    29442, 
    29445, 
    29448, 
    29451, 
    29454, 
    29457, 
    29460, 
    29463, 
    29466, 
    29469, 
    29472, 
    29475, 
    29478, 
    29481, 
    29484, 
    29487, 
    29490, 
    29493, 
    29496, 
    29499, 
    29502, 
    29505, 
    29508, 
    29511, 
    29514, 
    29517, 
    29520, 
    29523, 
    29526, 
    29529, 
    29532, 
    29535, 
    29538, 
    29541, 
    29544, 
    29547, 
    29550, 
    29553, 
    29556, 
    29559, 
    29562, 
    29565, 
    29568, 
    29571, 
    29574, 
    29577, 
    29580, 
    29583, 
    29586, 
    29589, 
    29592, 
    29595, 
    29598, 
    29601, 
    29604, 
    29607, 
    29610, 
    29613, 
    29616, 
    29619, 
    29622, 
    29625, 
    29628, 
    29631, 
    29634, 
    29637, 
    29640, 
    29643, 
    29646, 
    29649, 
    29652, 
    29655, 
    29658, 
    29661, 
    29664, 
    29667, 
    29670, 
    29673, 
    29676, 
    29679, 
    29682, 
    29685, 
    29688, 
    29691, 
    29694, 
    29697, 
    29700, 
    29703, 
    29706, 
    29709, 
    29712, 
    29715, 
    29718, 
    29721, 
    29724, 
    29727, 
    29730, 
    29733, 
    29736, 
    29739, 
    29742, 
    29745, 
    29748, 
    29751, 
    29754, 
    29757, 
    29760, 
    29763, 
    29766, 
    29769, 
    29772, 
    29775, 
    29778, 
    29781, 
    29784, 
    29787, 
    29790, 
    29793, 
    29796, 
    29799, 
    29802, 
    29805, 
    29808, 
    29811, 
    29814, 
    29817, 
    29820, 
    29823, 
    29826, 
    29829, 
    29832, 
    29835, 
    29838, 
    29841, 
    29844, 
    29847, 
    29850, 
    29853, 
    29856, 
    29859, 
    29862, 
    29865, 
    29868, 
    29871, 
    29874, 
    29877, 
    29880, 
    29883, 
    29886, 
    29889, 
    29892, 
    29895, 
    29898, 
    29901, 
    29904, 
    29907, 
    29910, 
    29913, 
    29916, 
    29919, 
    29922, 
    29925, 
    29928, 
    29931, 
    29934, 
    29937, 
    29940, 
    29943, 
    29946, 
    29949, 
    29952, 
    29955, 
    29958, 
    29961, 
    29964, 
    29967, 
    29970, 
    29973, 
    29976, 
    29979, 
    29982, 
    29985, 
    29988, 
    29991, 
    29994, 
    29997, 
    30000, 
    30003, 
    30006, 
    30009, 
    30012, 
    30015, 
    30018, 
    30021, 
    30024, 
    30027, 
    30030, 
    30033, 
    30036, 
    30039, 
    30042, 
    30045, 
    30048, 
    30051, 
    30054, 
    30057, 
    30060, 
    30063, 
    30066, 
    30069, 
    30072, 
    30075, 
    30078, 
    30081, 
    30084, 
    30087, 
    30090, 
    30093, 
    30096, 
    30099, 
    30102, 
    30105, 
    30108, 
    30111, 
    30114, 
    30117, 
    30120, 
    30123, 
    30126, 
    30129, 
    30132, 
    30135, 
    30138, 
    30141, 
    30144, 
    30147, 
    30150, 
    30153, 
    30156, 
    30159, 
    30162, 
    30165, 
    30168, 
    30171, 
    30174, 
    30177, 
    30180, 
    30183, 
    30186, 
    30189, 
    30192, 
    30195, 
    30198, 
    30201, 
    30204, 
    30207, 
    30210, 
    30213, 
    30216, 
    30219, 
    30222, 
    30225, 
    30228, 
    30231, 
    30234, 
    30237, 
    30240, 
    30243, 
    30246, 
    30249, 
    30252, 
    30255, 
    30258, 
    30261, 
    30264, 
    30267, 
    30270, 
    30273, 
    30276, 
    30279, 
    30282, 
    30285, 
    30288, 
    30291, 
    30294, 
    30297, 
    30300, 
    30303, 
    30306, 
    30309, 
    30312, 
    30315, 
    30318, 
    30321, 
    30324, 
    30327, 
    30330, 
    30333, 
    30336, 
    30339, 
    30342, 
    30345, 
    30348, 
    30351, 
    30354, 
    30357, 
    30360, 
    30363, 
    30366, 
    30369, 
    30372, 
    30375, 
    30378, 
    30381, 
    30384, 
    30387, 
    30390, 
    30393, 
    30396, 
    30399, 
    30402, 
    30405, 
    30408, 
    30411, 
    30414, 
    30417, 
    30420, 
    30423, 
    30426, 
    30429, 
    30432, 
    30435, 
    30438, 
    30441, 
    30444, 
    30447, 
    30450, 
    30453, 
    30456, 
    30459, 
    30462, 
    30465, 
    30468, 
    30471, 
    30474, 
    30477, 
    30480, 
    30483, 
    30486, 
    30489, 
    30492, 
    30495, 
    30498, 
    30501, 
    30504, 
    30507, 
    30510, 
    30513, 
    30516, 
    30519, 
    30522, 
    30525, 
    30528, 
    30531, 
    30534, 
    30537, 
    30540, 
    30543, 
    30546, 
    30549, 
    30552, 
    30555, 
    30558, 
    30561, 
    30564, 
    30567, 
    30570, 
    30573, 
    30576, 
    30579, 
    30582, 
    30585, 
    30588, 
    30591, 
    30594, 
    30597, 
    30600, 
    30603, 
    30606, 
    30609, 
    30612, 
    30615, 
    30618, 
    30621, 
    30624, 
    30627, 
    30630, 
    30633, 
    30636, 
    30639, 
    30642, 
    30645, 
    30648, 
    30651, 
    30654, 
    30657, 
    30660, 
    30663, 
    30666, 
    30669, 
    30672, 
    30675, 
    30678, 
    30681, 
    30684, 
    30687, 
    30690, 
    30693, 
    30696, 
    30699, 
    30702, 
    30705, 
    30708, 
    30711, 
    30714, 
    30717, 
    30720, 
    30723, 
    30726, 
    30729, 
    30732, 
    30735, 
    30738, 
    30741, 
    30744, 
    30747, 
    30750, 
    30753, 
    30756, 
    30759, 
    30762, 
    30765, 
    30768, 
    30771, 
    30774, 
    30777, 
    30780, 
    30783, 
    30786, 
    30789, 
    30792, 
    30795, 
    30798, 
    30801, 
    30804, 
    30807, 
    30810, 
    30813, 
    30816, 
    30819, 
    30822, 
    30825, 
    30828, 
    30831, 
    30834, 
    30837, 
    30840, 
    30843, 
    30846, 
    30849, 
    30852, 
    30855, 
    30858, 
    30861, 
    30864, 
    30867, 
    30870, 
    30873, 
    30876, 
    30879, 
    30882, 
    30885, 
    30888, 
    30891, 
    30894, 
    30897, 
    30900, 
    30903, 
    30906, 
    30909, 
    30912, 
    30915, 
    30918, 
    30921, 
    30924, 
    30927, 
    30930, 
    30933, 
    30936, 
    30939, 
    30942, 
    30945, 
    30948, 
    30951, 
    30954, 
    30957, 
    30960, 
    30963, 
    30966, 
    30969, 
    30972, 
    30975, 
    30978, 
    30981, 
    30984, 
    30987, 
    30990, 
    30993, 
    30996, 
    30999, 
    31002, 
    31005, 
    31008, 
    31011, 
    31014, 
    31017, 
    31020, 
    31023, 
    31026, 
    31029, 
    31032, 
    31035, 
    31038, 
    31041, 
    31044, 
    31047, 
    31050, 
    31053, 
    31056, 
    31059, 
    31062, 
    31065, 
    31068, 
    31071, 
    31074, 
    31077, 
    31080, 
    31083, 
    31086, 
    31089, 
    31092, 
    31095, 
    31098, 
    31101, 
    31104, 
    31107, 
    31110, 
    31113, 
    31116, 
    31119, 
    31122, 
    31125, 
    31128, 
    31131, 
    31134, 
    31137, 
    31140, 
    31143, 
    31146, 
    31149, 
    31152, 
    31155, 
    31158, 
    31161, 
    31164, 
    31167, 
    31170, 
    31173, 
    31176, 
    31179, 
    31182, 
    31185, 
    31188, 
    31191, 
    31194, 
    31197, 
    31200, 
    31203, 
    31206, 
    31209, 
    31212, 
    31215, 
    31218, 
    31221, 
    31224, 
    31227, 
    31230, 
    31233, 
    31236, 
    31239, 
    31242, 
    31245, 
    31248, 
    31251, 
    31254, 
    31257, 
    31260, 
    31263, 
    31266, 
    31269, 
    31272, 
    31275, 
    31278, 
    31281, 
    31284, 
    31287, 
    31290, 
    31293, 
    31296, 
    31299, 
    31302, 
    31305, 
    31308, 
    31311, 
    31314, 
    31317, 
    31320, 
    31323, 
    31326, 
    31329, 
    31332, 
    31335, 
    31338, 
    31341, 
    31344, 
    31347, 
    31350, 
    31353, 
    31356, 
    31359, 
    31362, 
    31365, 
    31368, 
    31371, 
    31374, 
    31377, 
    31380, 
    31383, 
    31386, 
    31389, 
    31392, 
    31395, 
    31398, 
    31401, 
    31404, 
    31407, 
    31410, 
    31413, 
    31416, 
    31419, 
    31422, 
    31425, 
    31428, 
    31431, 
    31434, 
    31437, 
    31440, 
    31443, 
    31446, 
    31449, 
    31452, 
    31455, 
    31458, 
    31461, 
    31464, 
    31467, 
    31470, 
    31473, 
    31476, 
    31479, 
    31482, 
    31485, 
    31488, 
    31491, 
    31494, 
    31497, 
    31500, 
    31503, 
    31506, 
    31509, 
    31512, 
    31515, 
    31518, 
    31521, 
    31524, 
    31527, 
    31530, 
    31533, 
    31536, 
    31539, 
    31542, 
    31545, 
    31548, 
    31551, 
    31554, 
    31557, 
    31560, 
    31563, 
    31566, 
    31569, 
    31572, 
    31575, 
    31578, 
    31581, 
    31584, 
    31587, 
    31590, 
    31593, 
    31596, 
    31599, 
    31602, 
    31605, 
    31608, 
    31611, 
    31614, 
    31617, 
    31620, 
    31623, 
    31626, 
    31629, 
    31632, 
    31635, 
    31638, 
    31641, 
    31644, 
    31647, 
    31650, 
    31653, 
    31656, 
    31659, 
    31662, 
    31665, 
    31668, 
    31671, 
    31674, 
    31677, 
    31680, 
    31683, 
    31686, 
    31689, 
    31692, 
    31695, 
    31698, 
    31701, 
    31704, 
    31707, 
    31710, 
    31713, 
    31716, 
    31719, 
    31722, 
    31725, 
    31728, 
    31731, 
    31734, 
    31737, 
    31740, 
    31743, 
    31746, 
    31749, 
    31752, 
    31755, 
    31758, 
    31761, 
    31764, 
    31767, 
    31770, 
    31773, 
    31776, 
    31779, 
    31782, 
    31785, 
    31788, 
    31791, 
    31794, 
    31797, 
    31800, 
    31803, 
    31806, 
    31809, 
    31812, 
    31815, 
    31818, 
    31821, 
    31824, 
    31827, 
    31830, 
    31833, 
    31836, 
    31839, 
    31842, 
    31845, 
    31848, 
    31851, 
    31854, 
    31857, 
    31860, 
    31863, 
    31866, 
    31869, 
    31872, 
    31875, 
    31878, 
    31881, 
    31884, 
    31887, 
    31890, 
    31893, 
    31896, 
    31899, 
    31902, 
    31905, 
    31908, 
    31911, 
    31914, 
    31917, 
    31920, 
    31923, 
    31926, 
    31929, 
    31932, 
    31935, 
    31938, 
    31941, 
    31944, 
    31947, 
    31950, 
    31953, 
    31956, 
    31959, 
    31962, 
    31965, 
    31968, 
    31971, 
    31974, 
    31977, 
    31980, 
    31983, 
    31986, 
    31989, 
    31992, 
    31995, 
    31998, 
    32001, 
    32004, 
    32007, 
    32010, 
    32013, 
    32016, 
    32019, 
    32022, 
    32025, 
    32028, 
    32031, 
    32034, 
    32037, 
    32040, 
    32043, 
    32046, 
    32049, 
    32052, 
    32055, 
    32058, 
    32061, 
    32064, 
    32067, 
    32070, 
    32073, 
    32076, 
    32079, 
    32082, 
    32085, 
    32088, 
    32091, 
    32094, 
    32097, 
    32100, 
    32103, 
    32106, 
    32109, 
    32112, 
    32115, 
    32118, 
    32121, 
    32124, 
    32127, 
    32130, 
    32133, 
    32136, 
    32139, 
    32142, 
    32145, 
    32148, 
    32151, 
    32154, 
    32157, 
    32160, 
    32163, 
    32166, 
    32169, 
    32172, 
    32175, 
    32178, 
    32181, 
    32184, 
    32187, 
    32190, 
    32193, 
    32196, 
    32199, 
    32202, 
    32205, 
    32208, 
    32211, 
    32214, 
    32217, 
    32220, 
    32223, 
    32226, 
    32229, 
    32232, 
    32235, 
    32238, 
    32241, 
    32244, 
    32247, 
    32250, 
    32253, 
    32256, 
    32259, 
    32262, 
    32265, 
    32268, 
    32271, 
    32274, 
    32277, 
    32280, 
    32283, 
    32286, 
    32289, 
    32292, 
    32295, 
    32298, 
    32301, 
    32304, 
    32307, 
    32310, 
    32313, 
    32316, 
    32319, 
    32322, 
    32325, 
    32328, 
    32331, 
    32334, 
    32337, 
    32340, 
    32343, 
    32346, 
    32349, 
    32352, 
    32355, 
    32358, 
    32361, 
    32364, 
    32367, 
    32370, 
    32373, 
    32376, 
    32379, 
    32382, 
    32385, 
    32388, 
    32391, 
    32394, 
    32397, 
    32400, 
    32403, 
    32406, 
    32409, 
    32412, 
    32415, 
    32418, 
    32421, 
    32424, 
    32427, 
    32430, 
    32433, 
    32436, 
    32439, 
    32442, 
    32445, 
    32448, 
    32451, 
    32454, 
    32457, 
    32460, 
    32463, 
    32466, 
    32469, 
    32472, 
    32475, 
    32478, 
    32481, 
    32484, 
    32487, 
    32490, 
    32493, 
    32496, 
    32499, 
    32502, 
    32505, 
    32508, 
    32511, 
    32514, 
    32517, 
    32520, 
    32523, 
    32526, 
    32529, 
    32532, 
    32535, 
    32538, 
    32541, 
    32544, 
    32547, 
    32550, 
    32553, 
    32556, 
    32559, 
    32562, 
    32565, 
    32568, 
    32571, 
    32574, 
    32577, 
    32580, 
    32583, 
    32586, 
    32589, 
    32592, 
    32595, 
    32598, 
    32601, 
    32604, 
    32607, 
    32610, 
    32613, 
    32616, 
    32619, 
    32622, 
    32625, 
    32628, 
    32631, 
    32634, 
    32637, 
    32640, 
    32643, 
    32646, 
    32649, 
    32652, 
    32655, 
    32658, 
    32661, 
    32664, 
    32667, 
    32670, 
    32673, 
    32676, 
    32679, 
    32682, 
    32685, 
    32688, 
    32691, 
    32694, 
    32697, 
    32700, 
    32703, 
    32706, 
    32709, 
    32712, 
    32715, 
    32718, 
    32721, 
    32724, 
    32727, 
    32730, 
    32733, 
    32736, 
    32739, 
    32742, 
    32745, 
    32748, 
    32751, 
    32754, 
    32757, 
    32760, 
    32763, 
    32766, 
    32769, 
    32772, 
    32775, 
    32778, 
    32781, 
    32784, 
    32787, 
    32790, 
    32793, 
    32796, 
    32799, 
    32802, 
    32805, 
    32808, 
    32811, 
    32814, 
    32817, 
    32820, 
    32823, 
    32826, 
    32829, 
    32832, 
    32835, 
    32838, 
    32841, 
    32844, 
    32847, 
    32850, 
    32853, 
    32856, 
    32859, 
    32862, 
    32865, 
    32868, 
    32871, 
    32874, 
    32877, 
    32880, 
    32883, 
    32886, 
    32889, 
    32892, 
    32895, 
    32898, 
    32901, 
    32904, 
    32907, 
    32910, 
    32913, 
    32916, 
    32919, 
    32922, 
    32925, 
    32928, 
    32931, 
    32934, 
    32937, 
    32940, 
    32943, 
    32946, 
    32949, 
    32952, 
    32955, 
    32958, 
    32961, 
    32964, 
    32967, 
    32970, 
    32973, 
    32976, 
    32979, 
    32982, 
    32985, 
    32988, 
    32991, 
    32994, 
    32997, 
    33000, 
    33003, 
    33006, 
    33009, 
    33012, 
    33015, 
    33018, 
    33021, 
    33024, 
    33027, 
    33030, 
    33033, 
    33036, 
    33039, 
    33042, 
    33045, 
    33048, 
    33051, 
    33054, 
    33057, 
    33060, 
    33063, 
    33066, 
    33069, 
    33072, 
    33075, 
    33078, 
    33081, 
    33084, 
    33087, 
    33090, 
    33093, 
    33096, 
    33099, 
    33102, 
    33105, 
    33108, 
    33111, 
    33114, 
    33117, 
    33120, 
    33123, 
    33126, 
    33129, 
    33132, 
    33135, 
    33138, 
    33141, 
    33144, 
    33147, 
    33150, 
    33153, 
    33156, 
    33159, 
    33162, 
    33165, 
    33168, 
    33171, 
    33174, 
    33177, 
    33180, 
    33183, 
    33186, 
    33189, 
    33192, 
    33195, 
    33198, 
    33201, 
    33204, 
    33207, 
    33210, 
    33213, 
    33216, 
    33219, 
    33222, 
    33225, 
    33228, 
    33231, 
    33234, 
    33237, 
    33240, 
    33243, 
    33246, 
    33249, 
    33252, 
    33255, 
    33258, 
    33261, 
    33264, 
    33267, 
    33270, 
    33273, 
    33276, 
    33279, 
    33282, 
    33285, 
    33288, 
    33291, 
    33294, 
    33297, 
    33300, 
    33303, 
    33306, 
    33309, 
    33312, 
    33315, 
    33318, 
    33321, 
    33324, 
    33327, 
    33330, 
    33333, 
    33336, 
    33339, 
    33342, 
    33345, 
    33348, 
    33351, 
    33354, 
    33357, 
    33360, 
    33363, 
    33366, 
    33369, 
    33372, 
    33375, 
    33378, 
    33381, 
    33384, 
    33387, 
    33390, 
    33393, 
    33396, 
    33399, 
    33402, 
    33405, 
    33408, 
    33411, 
    33414, 
    33417, 
    33420, 
    33423, 
    33426, 
    33429, 
    33432, 
    33435, 
    33438, 
    33441, 
    33444, 
    33447, 
    33450, 
    33453, 
    33456, 
    33459, 
    33462, 
    33465, 
    33468, 
    33471, 
    33474, 
    33477, 
    33480, 
    33483, 
    33486, 
    33489, 
    33492, 
    33495, 
    33498, 
    33501, 
    33504, 
    33507, 
    33510, 
    33513, 
    33516, 
    33519, 
    33522, 
    33525, 
    33528, 
    33531, 
    33534, 
    33537, 
    33540, 
    33543, 
    33546, 
    33549, 
    33552, 
    33555, 
    33558, 
    33561, 
    33564, 
    33567, 
    33570, 
    33573, 
    33576, 
    33579, 
    33582, 
    33585, 
    33588, 
    33591, 
    33594, 
    33597, 
    33600, 
    33603, 
    33606, 
    33609, 
    33612, 
    33615, 
    33618, 
    33621, 
    33624, 
    33627, 
    33630, 
    33633, 
    33636, 
    33639, 
    33642, 
    33645, 
    33648, 
    33651, 
    33654, 
    33657, 
    33660, 
    33663, 
    33666, 
    33669, 
    33672, 
    33675, 
    33678, 
    33681, 
    33684, 
    33687, 
    33690, 
    33693, 
    33696, 
    33699, 
    33702, 
    33705, 
    33708, 
    33711, 
    33714, 
    33717, 
    33720, 
    33723, 
    33726, 
    33729, 
    33732, 
    33735, 
    33738, 
    33741, 
    33744, 
    33747, 
    33750, 
    33753, 
    33756, 
    33759, 
    33762, 
    33765, 
    33768, 
    33771, 
    33774, 
    33777, 
    33780, 
    33783, 
    33786, 
    33789, 
    33792, 
    33795, 
    33798, 
    33801, 
    33804, 
    33807, 
    33810, 
    33813, 
    33816, 
    33819, 
    33822, 
    33825, 
    33828, 
    33831, 
    33834, 
    33837, 
    33840, 
    33843, 
    33846, 
    33849, 
    33852, 
    33855, 
    33858, 
    33861, 
    33864, 
    33867, 
    33870, 
    33873, 
    33876, 
    33879, 
    33882, 
    33885, 
    33888, 
    33891, 
    33894, 
    33897, 
    33900, 
    33903, 
    33906, 
    33909, 
    33912, 
    33915, 
    33918, 
    33921, 
    33924, 
    33927, 
    33930, 
    33933, 
    33936, 
    33939, 
    33942, 
    33945, 
    33948, 
    33951, 
    33954, 
    33957, 
    33960, 
    33963, 
    33966, 
    33969, 
    33972, 
    33975, 
    33978, 
    33981, 
    33984, 
    33987, 
    33990, 
    33993, 
    33996, 
    33999, 
    34002, 
    34005, 
    34008, 
    34011, 
    34014, 
    34017, 
    34020, 
    34023, 
    34026, 
    34029, 
    34032, 
    34035, 
    34038, 
    34041, 
    34044, 
    34047, 
    34050, 
    34053, 
    34056, 
    34059, 
    34062, 
    34065, 
    34068, 
    34071, 
    34074, 
    34077, 
    34080, 
    34083, 
    34086, 
    34089, 
    34092, 
    34095, 
    34098, 
    34101, 
    34104, 
    34107, 
    34110, 
    34113, 
    34116, 
    34119, 
    34122, 
    34125, 
    34128, 
    34131, 
    34134, 
    34137, 
    34140, 
    34143, 
    34146, 
    34149, 
    34152, 
    34155, 
    34158, 
    34161, 
    34164, 
    34167, 
    34170, 
    34173, 
    34176, 
    34179, 
    34182, 
    34185, 
    34188, 
    34191, 
    34194, 
    34197, 
    34200, 
    34203, 
    34206, 
    34209, 
    34212, 
    34215, 
    34218, 
    34221, 
    34224, 
    34227, 
    34230, 
    34233, 
    34236, 
    34239, 
    34242, 
    34245, 
    34248, 
    34251, 
    34254, 
    34257, 
    34260, 
    34263, 
    34266, 
    34269, 
    34272, 
    34275, 
    34278, 
    34281, 
    34284, 
    34287, 
    34290, 
    34293, 
    34296, 
    34299, 
    34302, 
    34305, 
    34308, 
    34311, 
    34314, 
    34317, 
    34320, 
    34323, 
    34326, 
    34329, 
    34332, 
    34335, 
    34338, 
    34341, 
    34344, 
    34347, 
    34350, 
    34353, 
    34356, 
    34359, 
    34362, 
    34365, 
    34368, 
    34371, 
    34374, 
    34377, 
    34380, 
    34383, 
    34386, 
    34389, 
    34392, 
    34395, 
    34398, 
    34401, 
    34404, 
    34407, 
    34410, 
    34413, 
    34416, 
    34419, 
    34422, 
    34425, 
    34428, 
    34431, 
    34434, 
    34437, 
    34440, 
    34443, 
    34446, 
    34449, 
    34452, 
    34455, 
    34458, 
    34461, 
    34464, 
    34467, 
    34470, 
    34473, 
    34476, 
    34479, 
    34482, 
    34485, 
    34488, 
    34491, 
    34494, 
    34497, 
    34500, 
    34503, 
    34506, 
    34509, 
    34512, 
    34515, 
    34518, 
    34521, 
    34524, 
    34527, 
    34530, 
    34533, 
    34536, 
    34539, 
    34542, 
    34545, 
    34548, 
    34551, 
    34554, 
    34557, 
    34560, 
    34563, 
    34566, 
    34569, 
    34572, 
    34575, 
    34578, 
    34581, 
    34584, 
    34587, 
    34590, 
    34593, 
    34596, 
    34599, 
    34602, 
    34605, 
    34608, 
    34611, 
    34614, 
    34617, 
    34620, 
    34623, 
    34626, 
    34629, 
    34632, 
    34635, 
    34638, 
    34641, 
    34644, 
    34647, 
    34650, 
    34653, 
    34656, 
    34659, 
    34662, 
    34665, 
    34668, 
    34671, 
    34674, 
    34677, 
    34680, 
    34683, 
    34686, 
    34689, 
    34692, 
    34695, 
    34698, 
    34701, 
    34704, 
    34707, 
    34710, 
    34713, 
    34716, 
    34719, 
    34722, 
    34725, 
    34728, 
    34731, 
    34734, 
    34737, 
    34740, 
    34743, 
    34746, 
    34749, 
    34752, 
    34755, 
    34758, 
    34761, 
    34764, 
    34767, 
    34770, 
    34773, 
    34776, 
    34779, 
    34782, 
    34785, 
    34788, 
    34791, 
    34794, 
    34797, 
    34800, 
    34803, 
    34806, 
    34809, 
    34812, 
    34815, 
    34818, 
    34821, 
    34824, 
    34827, 
    34830, 
    34833, 
    34836, 
    34839, 
    34842, 
    34845, 
    34848, 
    34851, 
    34854, 
    34857, 
    34860, 
    34863, 
    34866, 
    34869, 
    34872, 
    34875, 
    34878, 
    34881, 
    34884, 
    34887, 
    34890, 
    34893, 
    34896, 
    34899, 
    34902, 
    34905, 
    34908, 
    34911, 
    34914, 
    34917, 
    34920, 
    34923, 
    34926, 
    34929, 
    34932, 
    34935, 
    34938, 
    34941, 
    34944, 
    34947, 
    34950, 
    34953, 
    34956, 
    34959, 
    34962, 
    34965, 
    34968, 
    34971, 
    34974, 
    34977, 
    34980, 
    34983, 
    34986, 
    34989, 
    34992, 
    34995, 
    34998, 
    35001, 
    35004, 
    35007, 
    35010, 
    35013, 
    35016, 
    35019, 
    35022, 
    35025, 
    35028, 
    35031, 
    35034, 
    35037, 
    35040, 
    35043, 
    35046, 
    35049, 
    35052, 
    35055, 
    35058, 
    35061, 
    35064, 
    35067, 
    35070, 
    35073, 
    35076, 
    35079, 
    35082, 
    35085, 
    35088, 
    35091, 
    35094, 
    35097, 
    35100, 
    35103, 
    35106, 
    35109, 
    35112, 
    35115, 
    35118, 
    35121, 
    35124, 
    35127, 
    35130, 
    35133, 
    35136, 
    35139, 
    35142, 
    35145, 
    35148, 
    35151, 
    35154, 
    35157, 
    35160, 
    35163, 
    35166, 
    35169, 
    35172, 
    35175, 
    35178, 
    35181, 
    35184, 
    35187, 
    35190, 
    35193, 
    35196, 
    35199, 
    35202, 
    35205, 
    35208, 
    35211, 
    35214, 
    35217, 
    35220, 
    35223, 
    35226, 
    35229, 
    35232, 
    35235, 
    35238, 
    35241, 
    35244, 
    35247, 
    35250, 
    35253, 
    35256, 
    35259, 
    35262, 
    35265, 
    35268, 
    35271, 
    35274, 
    35277, 
    35280, 
    35283, 
    35286, 
    35289, 
    35292, 
    35295, 
    35298, 
    35301, 
    35304, 
    35307, 
    35310, 
    35313, 
    35316, 
    35319, 
    35322, 
    35325, 
    35328, 
    35331, 
    35334, 
    35337, 
    35340, 
    35343, 
    35346, 
    35349, 
    35352, 
    35355, 
    35358, 
    35361, 
    35364, 
    35367, 
    35370, 
    35373, 
    35376, 
    35379, 
    35382, 
    35385, 
    35388, 
    35391, 
    35394, 
    35397, 
    35400, 
    35403, 
    35406, 
    35409, 
    35412, 
    35415, 
    35418, 
    35421, 
    35424, 
    35427, 
    35430, 
    35433, 
    35436, 
    35439, 
    35442, 
    35445, 
    35448, 
    35451, 
    35454, 
    35457, 
    35460, 
    35463, 
    35466, 
    35469, 
    35472, 
    35475, 
    35478, 
    35481, 
    35484, 
    35487, 
    35490, 
    35493, 
    35496, 
    35499, 
    35502, 
    35505, 
    35508, 
    35511, 
    35514, 
    35517, 
    35520, 
    35523, 
    35526, 
    35529, 
    35532, 
    35535, 
    35538, 
    35541, 
    35544, 
    35547, 
    35550, 
    35553, 
    35556, 
    35559, 
    35562, 
    35565, 
    35568, 
    35571, 
    35574, 
    35577, 
    35580, 
    35583, 
    35586, 
    35589, 
    35592, 
    35595, 
    35598, 
    35601, 
    35604, 
    35607, 
    35610, 
    35613, 
    35616, 
    35619, 
    35622, 
    35625, 
    35628, 
    35631, 
    35634, 
    35637, 
    35640, 
    35643, 
    35646, 
    35649, 
    35652, 
    35655, 
    35658, 
    35661, 
    35664, 
    35667, 
    35670, 
    35673, 
    35676, 
    35679, 
    35682, 
    35685, 
    35688, 
    35691, 
    35694, 
    35697, 
    35700, 
    35703, 
    35706, 
    35709, 
    35712, 
    35715, 
    35718, 
    35721, 
    35724, 
    35727, 
    35730, 
    35733, 
    35736, 
    35739, 
    35742, 
    35745, 
    35748, 
    35751, 
    35754, 
    35757, 
    35760, 
    35763, 
    35766, 
    35769, 
    35772, 
    35775, 
    35778, 
    35781, 
    35784, 
    35787, 
    35790, 
    35793, 
    35796, 
    35799, 
    35802, 
    35805, 
    35808, 
    35811, 
    35814, 
    35817, 
    35820, 
    35823, 
    35826, 
    35829, 
    35832, 
    35835, 
    35838, 
    35841, 
    35844, 
    35847, 
    35850, 
    35853, 
    35856, 
    35859, 
    35862, 
    35865, 
    35868, 
    35871, 
    35874, 
    35877, 
    35880, 
    35883, 
    35886, 
    35889, 
    35892, 
    35895, 
    35898, 
    35901, 
    35904, 
    35907, 
    35910, 
    35913, 
    35916, 
    35919, 
    35922, 
    35925, 
    35928, 
    35931, 
    35934, 
    35937, 
    35940, 
    35943, 
    35946, 
    35949, 
    35952, 
    35955, 
    35958, 
    35961, 
    35964, 
    35967, 
    35970, 
    35973, 
    35976, 
    35979, 
    35982, 
    35985, 
    35988, 
    35991, 
    35994, 
    35997, 
    36000, 
    36003, 
    36006, 
    36009, 
    36012, 
    36015, 
    36018, 
    36021, 
    36024, 
    36027, 
    36030, 
    36033, 
    36036, 
    36039, 
    36042, 
    36045, 
    36048, 
    36051, 
    36054, 
    36057, 
    36060, 
    36063, 
    36066, 
    36069, 
    36072, 
    36075, 
    36078, 
    36081, 
    36084, 
    36087, 
    36090, 
    36093, 
    36096, 
    36099, 
    36102, 
    36105, 
    36108, 
    36111, 
    36114, 
    36117, 
    36120, 
    36123, 
    36126, 
    36129, 
    36132, 
    36135, 
    36138, 
    36141, 
    36144, 
    36147, 
    36150, 
    36153, 
    36156, 
    36159, 
    36162, 
    36165, 
    36168, 
    36171, 
    36174, 
    36177, 
    36180, 
    36183, 
    36186, 
    36189, 
    36192, 
    36195, 
    36198, 
    36201, 
    36204, 
    36207, 
    36210, 
    36213, 
    36216, 
    36219, 
    36222, 
    36225, 
    36228, 
    36231, 
    36234, 
    36237, 
    36240, 
    36243, 
    36246, 
    36249, 
    36252, 
    36255, 
    36258, 
    36261, 
    36264, 
    36267, 
    36270, 
    36273, 
    36276, 
    36279, 
    36282, 
    36285, 
    36288, 
    36291, 
    36294, 
    36297, 
    36300, 
    36303, 
    36306, 
    36309, 
    36312, 
    36315, 
    36318, 
    36321, 
    36324, 
    36327, 
    36330, 
    36333, 
    36336, 
    36339, 
    36342, 
    36345, 
    36348, 
    36351, 
    36354, 
    36357, 
    36360, 
    36363, 
    36366, 
    36369, 
    36372, 
    36375, 
    36378, 
    36381, 
    36384, 
    36387, 
    36390, 
    36393, 
    36396, 
    36399, 
    36402, 
    36405, 
    36408, 
    36411, 
    36414, 
    36417, 
    36420, 
    36423, 
    36426, 
    36429, 
    36432, 
    36435, 
    36438, 
    36441, 
    36444, 
    36447, 
    36450, 
    36453, 
    36456, 
    36459, 
    36462, 
    36465, 
    36468, 
    36471, 
    36474, 
    36477, 
    36480, 
    36483, 
    36486, 
    36489, 
    36492, 
    36495, 
    36498, 
    36501, 
    36504, 
    36507, 
    36510, 
    36513, 
    36516, 
    36519, 
    36522, 
    36525, 
    36528, 
    36531, 
    36534, 
    36537, 
    36540, 
    36543, 
    36546, 
    36549, 
    36552, 
    36555, 
    36558, 
    36561, 
    36564, 
    36567, 
    36570, 
    36573, 
    36576, 
    36579, 
    36582, 
    36585, 
    36588, 
    36591, 
    36594, 
    36597, 
    36600, 
    36603, 
    36606, 
    36609, 
    36612, 
    36615, 
    36618, 
    36621, 
    36624, 
    36627, 
    36630, 
    36633, 
    36636, 
    36639, 
    36642, 
    36645, 
    36648, 
    36651, 
    36654, 
    36657, 
    36660, 
    36663, 
    36666, 
    36669, 
    36672, 
    36675, 
    36678, 
    36681, 
    36684, 
    36687, 
    36690, 
    36693, 
    36696, 
    36699, 
    36702, 
    36705, 
    36708, 
    36711, 
    36714, 
    36717, 
    36720, 
    36723, 
    36726, 
    36729, 
    36732, 
    36735, 
    36738, 
    36741, 
    36744, 
    36747, 
    36750, 
    36753, 
    36756, 
    36759, 
    36762, 
    36765, 
    36768, 
    36771, 
    36774, 
    36777, 
    36780, 
    36783, 
    36786, 
    36789, 
    36792, 
    36795, 
    36798, 
    36801, 
    36804, 
    36807, 
    36810, 
    36813, 
    36816, 
    36819, 
    36822, 
    36825, 
    36828, 
    36831, 
    36834, 
    36837, 
    36840, 
    36843, 
    36846, 
    36849, 
    36852, 
    36855, 
    36858, 
    36861, 
    36864, 
    36867, 
    36870, 
    36873, 
    36876, 
    36879, 
    36882, 
    36885, 
    36888, 
    36891, 
    36894, 
    36897, 
    36900, 
    36903, 
    36906, 
    36909, 
    36912, 
    36915, 
    36918, 
    36921, 
    36924, 
    36927, 
    36930, 
    36933, 
    36936, 
    36939, 
    36942, 
    36945, 
    36948, 
    36951, 
    36954, 
    36957, 
    36960, 
    36963, 
    36966, 
    36969, 
    36972, 
    36975, 
    36978, 
    36981, 
    36984, 
    36987, 
    36990, 
    36993, 
    36996, 
    36999, 
    37002, 
    37005, 
    37008, 
    37011, 
    37014, 
    37017, 
    37020, 
    37023, 
    37026, 
    37029, 
    37032, 
    37035, 
    37038, 
    37041, 
    37044, 
    37047, 
    37050, 
    37053, 
    37056, 
    37059, 
    37062, 
    37065, 
    37068, 
    37071, 
    37074, 
    37077, 
    37080, 
    37083, 
    37086, 
    37089, 
    37092, 
    37095, 
    37098, 
    37101, 
    37104, 
    37107, 
    37110, 
    37113, 
    37116, 
    37119, 
    37122, 
    37125, 
    37128, 
    37131, 
    37134, 
    37137, 
    37140, 
    37143, 
    37146, 
    37149, 
    37152, 
    37155, 
    37158, 
    37161, 
    37164, 
    37167, 
    37170, 
    37173, 
    37176, 
    37179, 
    37182, 
    37185, 
    37188, 
    37191, 
    37194, 
    37197, 
    37200, 
    37203, 
    37206, 
    37209, 
    37212, 
    37215, 
    37218, 
    37221, 
    37224, 
    37227, 
    37230, 
    37233, 
    37236, 
    37239, 
    37242, 
    37245, 
    37248, 
    37251, 
    37254, 
    37257, 
    37260, 
    37263, 
    37266, 
    37269, 
    37272, 
    37275, 
    37278, 
    37281, 
    37284, 
    37287, 
    37290, 
    37293, 
    37296, 
    37299, 
    37302, 
    37305, 
    37308, 
    37311, 
    37314, 
    37317, 
    37320, 
    37323, 
    37326, 
    37329, 
    37332, 
    37335, 
    37338, 
    37341, 
    37344, 
    37347, 
    37350, 
    37353, 
    37356, 
    37359, 
    37362, 
    37365, 
    37368, 
    37371, 
    37374, 
    37377, 
    37380, 
    37383, 
    37386, 
    37389, 
    37392, 
    37395, 
    37398, 
    37401, 
    37404, 
    37407, 
    37410, 
    37413, 
    37416, 
    37419, 
    37422, 
    37425, 
    37428, 
    37431, 
    37434, 
    37437, 
    37440, 
    37443, 
    37446, 
    37449, 
    37452, 
    37455, 
    37458, 
    37461, 
    37464, 
    37467, 
    37470, 
    37473, 
    37476, 
    37479, 
    37482, 
    37485, 
    37488, 
    37491, 
    37494, 
    37497, 
    37500, 
    37503, 
    37506, 
    37509, 
    37512, 
    37515, 
    37518, 
    37521, 
    37524, 
    37527, 
    37530, 
    37533, 
    37536, 
    37539, 
    37542, 
    37545, 
    37548, 
    37551, 
    37554, 
    37557, 
    37560, 
    37563, 
    37566, 
    37569, 
    37572, 
    37575, 
    37578, 
    37581, 
    37584, 
    37587, 
    37590, 
    37593, 
    37596, 
    37599, 
    37602, 
    37605, 
    37608, 
    37611, 
    37614, 
    37617, 
    37620, 
    37623, 
    37626, 
    37629, 
    37632, 
    37635, 
    37638, 
    37641, 
    37644, 
    37647, 
    37650, 
    37653, 
    37656, 
    37659, 
    37662, 
    37665, 
    37668, 
    37671, 
    37674, 
    37677, 
    37680, 
    37683, 
    37686, 
    37689, 
    37692, 
    37695, 
    37698, 
    37701, 
    37704, 
    37707, 
    37710, 
    37713, 
    37716, 
    37719, 
    37722, 
    37725, 
    37728, 
    37731, 
    37734, 
    37737, 
    37740, 
    37743, 
    37746, 
    37749, 
    37752, 
    37755, 
    37758, 
    37761, 
    37764, 
    37767, 
    37770, 
    37773, 
    37776, 
    37779, 
    37782, 
    37785, 
    37788, 
    37791, 
    37794, 
    37797, 
    37800, 
    37803, 
    37806, 
    37809, 
    37812, 
    37815, 
    37818, 
    37821, 
    37824, 
    37827, 
    37830, 
    37833, 
    37836, 
    37839, 
    37842, 
    37845, 
    37848, 
    37851, 
    37854, 
    37857, 
    37860, 
    37863, 
    37866, 
    37869, 
    37872, 
    37875, 
    37878, 
    37881, 
    37884, 
    37887, 
    37890, 
    37893, 
    37896, 
    37899, 
    37902, 
    37905, 
    37908, 
    37911, 
    37914, 
    37917, 
    37920, 
    37923, 
    37926, 
    37929, 
    37932, 
    37935, 
    37938, 
    37941, 
    37944, 
    37947, 
    37950, 
    37953, 
    37956, 
    37959, 
    37962, 
    37965, 
    37968, 
    37971, 
    37974, 
    37977, 
    37980, 
    37983, 
    37986, 
    37989, 
    37992, 
    37995, 
    37998, 
    38001, 
    38004, 
    38007, 
    38010, 
    38013, 
    38016, 
    38019, 
    38022, 
    38025, 
    38028, 
    38031, 
    38034, 
    38037, 
    38040, 
    38043, 
    38046, 
    38049, 
    38052, 
    38055, 
    38058, 
    38061, 
    38064, 
    38067, 
    38070, 
    38073, 
    38076, 
    38079, 
    38082, 
    38085, 
    38088, 
    38091, 
    38094, 
    38097, 
    38100, 
    38103, 
    38106, 
    38109, 
    38112, 
    38115, 
    38118, 
    38121, 
    38124, 
    38127, 
    38130, 
    38133, 
    38136, 
    38139, 
    38142, 
    38145, 
    38148, 
    38151, 
    38154, 
    38157, 
    38160, 
    38163, 
    38166, 
    38169, 
    38172, 
    38175, 
    38178, 
    38181, 
    38184, 
    38187, 
    38190, 
    38193, 
    38196, 
    38199, 
    38202, 
    38205, 
    38208, 
    38211, 
    38214, 
    38217, 
    38220, 
    38223, 
    38226, 
    38229, 
    38232, 
    38235, 
    38238, 
    38241, 
    38244, 
    38247, 
    38250, 
    38253 ;

 vertices.elevation = 
    780.780549531285, 
    1532.01409571516, 
    1170.62423732871, 
    1245.47898421317, 
    1386.17110983712, 
    1413.63980032655, 
    849.169647067285, 
    468.687296639813, 
    154.119670098759, 
    169.531916979818, 
    622.178889792443, 
    1202.59120153363, 
    1024.74734731558, 
    363.352368334566, 
    1433.88415832497, 
    1286.70089410275, 
    1719.42589559484, 
    1500.51557650079, 
    797.304238643797, 
    590.906971769848, 
    546.199408348328, 
    172.191147081167, 
    782.977420691792, 
    1154.10344339783, 
    139.191096070685, 
    1222.22960860587, 
    1445.81036706738, 
    1925.68525330069, 
    1754.48404124345, 
    1952.98926916511, 
    1410.19601680461, 
    1227.77145411519, 
    1133.42936630709, 
    1683.41203363333, 
    1141.21714290294, 
    1688.27301381235, 
    2158.57213717519, 
    1376.21413125465, 
    2103.45826886044, 
    0, 
    1225.63132112663, 
    1598.01754273982, 
    1253.16242690395, 
    1159.47435103054, 
    1196.17174813576, 
    1120.57777639485, 
    473.294465934207, 
    1020.01310325975, 
    1121.18123848938, 
    476.461925330178, 
    1304.89825627146, 
    2114.71290456493, 
    1768.9370217013, 
    1668.00787389144, 
    2002.40863742691, 
    972.76184341989, 
    1289.55670870708, 
    1754.43493007791, 
    2098.3260835934, 
    1431.70829820573, 
    1793.73368227324, 
    1456.1539570058, 
    771.765834601108, 
    57.6882343592817, 
    786.532963319033, 
    1165.25629528622, 
    638.761175835182, 
    1330.75022175135, 
    1198.09720390356, 
    635.057855244825, 
    394.860730810034, 
    1504.74120233327, 
    553.886290510005, 
    1598.78037156449, 
    1299.36982325373, 
    1180.5206792935, 
    130.707444152233, 
    1008.48484451861, 
    607.314141260553, 
    1249.56391026339, 
    1416.89997866737, 
    1636.8867191291, 
    437.655578557772, 
    795.502144461487, 
    1723.07214442483, 
    1586.57570796782, 
    840.048853344145, 
    300.310465126073, 
    219.658594440977, 
    1108.64604265551, 
    1631.87650156752, 
    1559.95603626508, 
    100.354566292252, 
    1221.05779119065, 
    1669.30978707094, 
    1468.18752794046, 
    959.970981463065, 
    891.969580863522, 
    987.602774939156, 
    364.949192956448, 
    0.103616813294233, 
    1245.70253377693, 
    757.674717626615, 
    613.690048590083, 
    861.470584583383, 
    256.355901959157, 
    735.953367511202, 
    507.213621592659, 
    450.747937936396, 
    624.126863425438, 
    584.085487606264, 
    1037.91889073778, 
    182.081879433114, 
    711.322926326283, 
    0, 
    1247.52317195965, 
    2091.28597160946, 
    653.279661553732, 
    490.804752420833, 
    2066.4120682014, 
    1206.14562894125, 
    907.122733467442, 
    136.931510417998, 
    721.984973301164, 
    1613.82183357273, 
    1710.04377221856, 
    1429.18254661434, 
    12.3653043151311, 
    723.869036085399, 
    1057.92246336517, 
    509.743930573189, 
    1144.59910504791, 
    483.293750051355, 
    1026.30789804339, 
    1460.94774701901, 
    1279.41625309963, 
    1792.10715948972, 
    539.017009504076, 
    656.139924541979, 
    112.34065683351, 
    1158.83294985126, 
    902.746721097106, 
    338.022575428407, 
    123.303703198628, 
    89.7797604305507, 
    0.103616813294233, 
    412.450622920113, 
    333.824906665075, 
    20.1763072416012, 
    0.103616813294233, 
    1236.34861061607, 
    472.410335911589, 
    647.695524788355, 
    326.778561068197, 
    1039.71944036181, 
    455.961108037561, 
    0.103616813294233, 
    952.964919620454, 
    902.92458081571, 
    1374.90772786696, 
    281.983151859866, 
    367.653297603889, 
    718.32519707952, 
    191.790087285549, 
    812.069366185414, 
    1052.95921179332, 
    343.369318697449, 
    771.24145216217, 
    226.588162818895, 
    899.433439122673, 
    871.752226698494, 
    737.552192342701, 
    724.33025470882, 
    124.675963197266, 
    735.914778039291, 
    627.430804602942, 
    59.2595992943223, 
    499.624700665787, 
    101.21242236166, 
    301.077656808106, 
    486.261293536691, 
    437.16564252137, 
    251.989503817311, 
    0.16585904238136, 
    446.18513317174, 
    248.623584743531, 
    174.303488135033, 
    0, 
    462.973983900036, 
    0, 
    80.8468962840409, 
    0.103616813294233, 
    205.862568742801, 
    212.068585114503, 
    134.01618863388, 
    0.943289424530187, 
    0, 
    293.994918765746, 
    172.934428981064, 
    884.592873314219, 
    594.319484895399, 
    1511.19848281819, 
    759.780840719335, 
    523.287235165142, 
    853.188210969359, 
    1581.72820509131, 
    790.706819716267, 
    874.76832300374, 
    968.672949967565, 
    0, 
    682.946283105009, 
    308.456010532437, 
    691.901635821519, 
    1153.26352964347, 
    5.65663892473168, 
    311.059041657405, 
    424.873415148969, 
    316.914146357566, 
    447.590356762132, 
    0, 
    258.422543630154, 
    44.5238510414212, 
    475.92802665821, 
    408.969770281493, 
    979.727478573501, 
    330.927998372397, 
    250.834668051122, 
    407.084366735336, 
    413.968094478888, 
    924.088434840224, 
    1299.54610811637, 
    1606.18540833027, 
    305.330843301895, 
    560.797026054183, 
    807.525053364174, 
    1613.0939240412, 
    1399.04171342759, 
    1673.91533102934, 
    976.163105602816, 
    1685.3635621734, 
    1257.56910347233, 
    339.177500194798, 
    187.666259382345, 
    1244.52290595398, 
    1492.07550501372, 
    433.861098773297, 
    1303.9107599553, 
    1581.64228933605, 
    707.030525354782, 
    1063.66215528424, 
    435.104229570397, 
    390.730972719743, 
    237.327842660971, 
    94.2023291370126, 
    455.355433101879, 
    463.130709803414, 
    51.9686012703483, 
    329.717194644408, 
    887.075221879567, 
    923.765427438207, 
    1120.75207228138, 
    745.551973102166, 
    624.374176893016, 
    812.548144497132, 
    832.050114248601, 
    491.945325023326, 
    741.064888226767, 
    861.920972631109, 
    845.951741229952, 
    691.970607634867, 
    714.854662320884, 
    599.269192879554, 
    235.966975529286, 
    255.126760022794, 
    899.888832512899, 
    1017.78168472146, 
    309.24320517106, 
    1610.15510923542, 
    792.904645583921, 
    1324.44493569494, 
    972.267730594091, 
    563.389677916017, 
    1175.84650492411, 
    229.406753799276, 
    525.373778763055, 
    1082.72377114318, 
    1071.19259885633, 
    1114.9268481104, 
    851.92674213185, 
    420.315868241836, 
    875.795679989486, 
    71.30801143352, 
    900.260371406044, 
    958.58383026407, 
    522.756756505366, 
    901.125296192609, 
    817.364327932235, 
    849.086914938815, 
    1211.05451680004, 
    651.664252622987, 
    311.701603065974, 
    705.974424845059, 
    629.740674951714, 
    966.690562365651, 
    482.962619168652, 
    228.245854356948, 
    816.836947279219, 
    831.976015279309, 
    1011.17911563126, 
    722.096698383452, 
    742.086405356043, 
    380.140730602557, 
    459.07338671748, 
    619.347160866558, 
    583.753526868828, 
    603.81883111349, 
    355.860773100211, 
    525.517288599275, 
    234.166227203615, 
    156.025284135283, 
    413.477460669015, 
    256.095355691675, 
    442.68761259559, 
    328.308017786826, 
    248.818669333184, 
    511.449258977676, 
    476.890257891872, 
    481.731228669425, 
    99.196499136528, 
    372.996180277824, 
    452.621436403766, 
    672.031651815386, 
    612.082885432841, 
    632.371937387418, 
    655.348535549755, 
    804.645433808095, 
    862.198446510862, 
    696.344714571092, 
    0.103616813294233, 
    1660.75670878575, 
    806.434838293984, 
    1889.64743630912, 
    1815.77330568645, 
    385.337774940322, 
    1676.18672434451, 
    1619.28442230725, 
    303.560578904281, 
    608.807194627692, 
    1667.71729597719, 
    1127.24809896275, 
    1367.78310335039, 
    494.9666947345, 
    0.103616813294233, 
    26.7786836015193, 
    0.103616813294233, 
    275.299082089045, 
    315.245179172755, 
    551.147048405711, 
    140.66842285589, 
    59.3701269392051, 
    462.700574065009, 
    0.103616813294233, 
    37.1353012801088, 
    290.598117041338, 
    0.103616813294233, 
    91.3921783052576, 
    404.441205657696, 
    0.103616813294233, 
    0, 
    28.3802275366551, 
    769.904573606227, 
    928.140074309448, 
    0.103616813294233, 
    209.538162929116, 
    0.198235565538615, 
    0.103616813294233, 
    158.369636645289, 
    0, 
    0.103616813294233, 
    385.444048368876, 
    543.967734635597, 
    142.459649945802, 
    200.193978235062, 
    455.639799922203, 
    43.5964293699801, 
    818.879920363285, 
    0.103616813294233, 
    184.916120878721, 
    27.8424040245806, 
    3.37158348095868, 
    37.2247087809381, 
    231.70517634087, 
    542.15605459022, 
    0.114146319770051, 
    0, 
    22.1033874692085, 
    150.025603665265, 
    37.2277240814259, 
    630.373080293902, 
    406.673960924493, 
    33.1176855739957, 
    361.121765104557, 
    415.98964487002, 
    507.695812576516, 
    643.152014235606, 
    410.610267169818, 
    658.368288588738, 
    284.11867335006, 
    814.300556794173, 
    56.7051469245636, 
    555.296807970423, 
    171.474258377023, 
    640.5314999576, 
    186.594515737337, 
    255.21753843251, 
    659.94549325924, 
    358.430810789662, 
    739.675965175397, 
    51.2342090600183, 
    279.492239379966, 
    0, 
    393.033639157233, 
    9.77118418817944, 
    123.938291180019, 
    200.217865696829, 
    724.777064695603, 
    610.296517034418, 
    662.631185993868, 
    661.482264659053, 
    816.612831581813, 
    594.136758172744, 
    732.318176640923, 
    601.778827806273, 
    560.377161475101, 
    263.711392161181, 
    0.103616813294233, 
    34.7850004775829, 
    71.980064390531, 
    56.1821707658575, 
    516.29102354405, 
    232.246281761409, 
    453.450033966655, 
    791.896765551912, 
    707.718738716851, 
    754.553044335244, 
    245.499522698673, 
    219.145253318826, 
    224.478894695625, 
    75.7013159248113, 
    704.005382568001, 
    871.053515494206, 
    19.7941968099967, 
    874.571657624422, 
    558.592619535944, 
    942.870688683035, 
    687.345555227799, 
    989.492867422466, 
    1012.94419793172, 
    688.470853982506, 
    237.612687741817, 
    491.519817438758, 
    802.819150944781, 
    293.462520272007, 
    710.406398115239, 
    792.582506773954, 
    723.378603644292, 
    614.202168847804, 
    304.75975403674, 
    965.103379353291, 
    29.3939507029726, 
    630.031517367665, 
    200.672666433166, 
    591.896787584681, 
    802.985708522517, 
    494.111978393806, 
    587.328040559763, 
    46.7357787632238, 
    34.8431994376753, 
    720.656243151442, 
    121.924233502235, 
    22.5447759439748, 
    281.27368912392, 
    840.254399092132, 
    770.74469333423, 
    546.898965911615, 
    647.181477367708, 
    766.529790980823, 
    443.558714382461, 
    38.9456149116516, 
    584.978617849408, 
    1024.93413818513, 
    364.759078652802, 
    1090.33239354867, 
    941.759208930037, 
    1026.17305853466, 
    297.601463434036, 
    858.133180875932, 
    798.972873757161, 
    801.667063150944, 
    161.445611354183, 
    728.557287790379, 
    926.143764243146, 
    950.600452224872, 
    531.916731755676, 
    41.2901623264582, 
    813.574948318623, 
    652.028131105114, 
    610.990644145841, 
    225.904125827038, 
    301.124934069379, 
    605.003444688816, 
    921.060616584301, 
    455.527286134963, 
    913.61966867044, 
    893.753701557331, 
    870.528102563568, 
    755.72725030148, 
    606.507414679754, 
    372.852710888715, 
    776.113829256583, 
    271.388749709073, 
    418.433612589703, 
    569.324170250964, 
    678.165960650713, 
    531.478014067028, 
    250.904915781765, 
    160.221041752295, 
    675.951367671008, 
    0.184402342630044, 
    905.750839797864, 
    33.4760884788146, 
    33.2974846607244, 
    760.716064856385, 
    109.135364243612, 
    155.208858687676, 
    82.3345651081697, 
    505.38775780235, 
    0.103616813294233, 
    0.103616813294233, 
    270.410860739704, 
    29.2050978844217, 
    154.310784628847, 
    372.36980882043, 
    601.62173723822, 
    84.0781187577275, 
    405.998567223335, 
    332.341049695539, 
    425.411885361883, 
    413.940739134842, 
    483.333133619282, 
    144.41980246846, 
    187.513626660277, 
    145.943096511313, 
    117.859640555155, 
    0.103616813294233, 
    78.8846134598648, 
    244.066249828057, 
    655.142586246658, 
    326.878750529057, 
    716.472102262312, 
    1343.06015794721, 
    1289.21765575424, 
    1176.44210258476, 
    1556.90068757014, 
    770.061100284977, 
    877.451381770738, 
    363.238808107918, 
    1176.83851345201, 
    1239.47600232319, 
    1236.00454205236, 
    2001.92938641893, 
    1506.59963407655, 
    1413.00417411666, 
    1500.85535813224, 
    1552.93501508053, 
    869.982527781452, 
    667.25298360667, 
    386.475644914394, 
    77.4018090388008, 
    374.91880519427, 
    681.935908543667, 
    895.18691048827, 
    392.893631450758, 
    813.284308945824, 
    1144.78909751734, 
    1209.19328669866, 
    1482.9493005011, 
    876.274418668234, 
    1106.41357885668, 
    569.897946645775, 
    1096.17234601136, 
    897.937595140184, 
    692.251542568624, 
    1345.36920038445, 
    843.616377518161, 
    1240.71395247031, 
    1097.19268269094, 
    679.475003566603, 
    1311.667499778, 
    1018.65026404223, 
    1528.2724520079, 
    657.074118328677, 
    581.656957524668, 
    126.023052914822, 
    712.017143214851, 
    1547.61414862089, 
    1730.50152983241, 
    573.842368222948, 
    411.075844390855, 
    224.939871880797, 
    954.193335346523, 
    891.893699027945, 
    755.677788562589, 
    171.509491716333, 
    553.03432745804, 
    790.183703388623, 
    951.849699521608, 
    736.287761072493, 
    639.477885438403, 
    620.332535838878, 
    1385.83773920523, 
    741, 
    833.991919534343, 
    916.39973530665, 
    733.855983059964, 
    600.540609354131, 
    600.638121452454, 
    433.818842112698, 
    399.452206331065, 
    164.82224511514, 
    492.432538729508, 
    506.939091202746, 
    72.3348489350441, 
    1346.00209124732, 
    1655.23781214374, 
    633.327518587617, 
    418.691716803688, 
    438.248566420356, 
    0.103616813294233, 
    0.172631996554792, 
    205.813522443366, 
    858.41854017801, 
    664.650081317738, 
    59.3530296270286, 
    58.4603273656651, 
    306.867458143404, 
    356.96973579017, 
    1096.90069022819, 
    36.3969504109504, 
    830.808344156255, 
    241.555614725533, 
    489.183342961932, 
    245.707644758878, 
    488.989132814193, 
    0.103616813294233, 
    423.582571009177, 
    123.155098026606, 
    70.9303235785266, 
    140.540159759145, 
    1057.88240673869, 
    1071.54733861258, 
    474.328808686331, 
    1019.34672878744, 
    936.993340118166, 
    2613.20950797002, 
    1169.50606087838, 
    986.761068583899, 
    1612.40195540329, 
    985.045768983241, 
    2633, 
    1175.18420938958, 
    2319.70269207277, 
    2199.61710763486, 
    1185.50280167524, 
    2107.7065646472, 
    2780.23087662805, 
    2867, 
    2091.15637554926, 
    26.6818260315372, 
    2482, 
    680.34048297429, 
    1690.45368365199, 
    2678.57984405199, 
    2279.0668104982, 
    2016.63868044437, 
    864.869781055077, 
    468.42995866602, 
    2283.90642857467, 
    3126.94681476455, 
    2324.44442418258, 
    1273.70055239499, 
    2552.41636632694, 
    3017.44981952453, 
    2606.73572919621, 
    2147.4276086969, 
    1129.61989317342, 
    969.625867509347, 
    1793.98957853888, 
    2057, 
    2788.59338686784, 
    1235.40414067986, 
    804.212443737405, 
    1420.72467964249, 
    698.242290696862, 
    683.530747820741, 
    2754.09922017784, 
    1455.5720035458, 
    3190, 
    2409.29282580101, 
    1361.59192352667, 
    2171.66773150859, 
    2153.18192721447, 
    1690.88011936642, 
    2031.44005097254, 
    2041.57484956469, 
    1935.51322300145, 
    2635.51994384995, 
    867.565837753083, 
    2134.96564730701, 
    2129.66535513179, 
    1609.57167159174, 
    831.636245603136, 
    2906, 
    2985.351305432, 
    2358.06144439846, 
    1483.87465846803, 
    2709, 
    3091, 
    1007.65986795797, 
    2061.68897179048, 
    2183.74837674919, 
    2301.05565807281, 
    2482.30246268869, 
    1606.14644446906, 
    2186, 
    2638, 
    958.492834840789, 
    2296.43506673184, 
    2171.9991001022, 
    1670.02102065054, 
    1114.04676696323, 
    1225.93489616787, 
    2910.00041105024, 
    2244.54017319862, 
    2439.73621423217, 
    2642.48549590781, 
    1898.78030144277, 
    2691.00062220395, 
    2002.86981852829, 
    2844, 
    1937.5229431577, 
    2778.50550488586, 
    1020.81339531791, 
    2426.172199003, 
    1010.44893567904, 
    2337.94897602102, 
    2082, 
    1329.08818122782, 
    2988.82816705284, 
    3109, 
    2281.2529614943, 
    3187, 
    2632.17344958879, 
    2603, 
    3217.06926507729, 
    1210.87859239053, 
    1253.95184019684, 
    2150.43595105867, 
    1033.68129099915, 
    2877, 
    1659.168812153, 
    1901.65335499669, 
    2174.02016536684, 
    903.867250581267, 
    1415.77503859801, 
    2881, 
    3061, 
    1312.19223664719, 
    1437.22226588866, 
    2526.15516400522, 
    2477.48014410121, 
    1578.82767939682, 
    2808.77630379082, 
    1093.53380173324, 
    1959.22032000307, 
    2045.27255080531, 
    1834.55555284548, 
    1335.30777809587, 
    1927.03276407737, 
    2855.95571555217, 
    1689.75468272428, 
    629.045603486395, 
    1998.58165922175, 
    2752.70344314287, 
    2447.67980915638, 
    1403.67030601546, 
    1803.78401080959, 
    3065, 
    1208.45873991924, 
    1284.92897063977, 
    1342.00490975146, 
    1608.47602683317, 
    1897.22601163802, 
    1482.37508540966, 
    3020.27233788272, 
    2829.72108121672, 
    2723, 
    1734, 
    1585.92250364647, 
    690.660214253954, 
    2635.04124511539, 
    546.680947423841, 
    1218.42654531699, 
    1703.69117486504, 
    2541.21569989269, 
    3155, 
    2413.33832496526, 
    1746.28854723964, 
    2887, 
    652.296174350174, 
    2657.49026644321, 
    2453.76553609269, 
    1542.53005918951, 
    1971.74915576521, 
    2084.01764313584, 
    2172.75784459637, 
    2642.31583099955, 
    1037.23778453536, 
    1744.72381535781, 
    2993, 
    736.853571662719, 
    1009.79259188693, 
    1350.03092225152, 
    1587.50256969185, 
    1858.74765000257, 
    374.575430548122, 
    2432, 
    2097.9143855154, 
    1503.01832883452, 
    1562, 
    1492.44328198405, 
    1995, 
    1627.35574498682, 
    3169, 
    2323.43852467568, 
    1913.03931175476, 
    1421.79461962361, 
    2854.55435566818, 
    1869.02471289576, 
    2508.02940519795, 
    1153.31272088992, 
    2697.50998280574, 
    1937.7773395503, 
    794.681329392749, 
    1763.98982820033, 
    2007.03766561058, 
    1435.21772648049, 
    1912.92901181807, 
    1515.62345908466, 
    3243, 
    1012.25546820399, 
    2924.02363226085, 
    1770.36052283627, 
    1929.54472147928, 
    2399.47466950074, 
    2049.02373735279, 
    1510.11960059217, 
    2421.52982546255, 
    1758.77438083738, 
    2521.70686142359, 
    1009.14706003093, 
    2887.68676796812, 
    2365.76566783122, 
    1239.93655117875, 
    942.702271221521, 
    912.484015687818, 
    2360, 
    1823.68120792876, 
    2585, 
    2216.06649687456, 
    1746.92023221208, 
    489.238696575746, 
    1684.63504316341, 
    2283.34320530837, 
    1942.1237192582, 
    2150.98734866636, 
    930.183186868963, 
    2121.89928311094, 
    2058.08743308694, 
    1695.08707384304, 
    1833.66528480347, 
    2450, 
    3140, 
    1607.26188995621, 
    2798.60515449358, 
    2820.13048832319, 
    577.926655178915, 
    2352.95181409757, 
    2513, 
    1973.57645287891, 
    1512.8244162358, 
    887.059794236915, 
    1726.15621252903, 
    835.275106303254, 
    1435.84597953469, 
    488.239064340547, 
    1318.01503113908, 
    843.218988242524, 
    577.407095484354, 
    2266.61217271004, 
    1476.36096220967, 
    3154.30706285748, 
    1801.13179376099, 
    2475.57726918902, 
    2532.02013852372, 
    2396, 
    986.929539334794, 
    1817.89587015727, 
    2758.1199629305, 
    237.706066132661, 
    2709.98340193074, 
    2020.55939016812, 
    2076, 
    1305.43849351619, 
    2995, 
    3182, 
    1786.26581614864, 
    1284.64088527704, 
    2832.44465715722, 
    2799, 
    2943.47949362854, 
    1924.64614240276, 
    1379.16029441087, 
    2464.05310880521, 
    1921.37054129704, 
    1632, 
    2888, 
    1500.18127175636, 
    2487.88525081733, 
    1984.44097659075, 
    1413.12847045621, 
    1172.93131739554, 
    2600, 
    2747.23666395398, 
    2192.00693881258, 
    2029.07101181115, 
    2450.0936289388, 
    2991.95452229469, 
    2137.49322435043, 
    729.413103627573, 
    2566.00090914637, 
    1583.48212894861, 
    1122.69376805171, 
    1924.83855083784, 
    35.5992338967595, 
    1935.11693883648, 
    2763.44336499101, 
    3009, 
    2926, 
    1059.232906121, 
    2553.02687337406, 
    3205, 
    690.419141241487, 
    523.913941170317, 
    2359, 
    2235.15057538105, 
    1887.6606443068, 
    1636.14265541923, 
    2679.09466279069, 
    1032.56131153147, 
    1908.38439340148, 
    2176.95106644133, 
    1293.17919789094, 
    2343, 
    1259.17376584433, 
    1223.72942853752, 
    630.720344218053, 
    2813.83295490082, 
    3165, 
    49.3053423472021, 
    1642.24502056231, 
    1619.71833860781, 
    1824.59083120188, 
    1267.05824676468, 
    1530.26406691713, 
    2060, 
    1872.87551594768, 
    1603.25931608244, 
    2925.15234519778, 
    1684.55834816343, 
    1414.92140075415, 
    2465.29724367329, 
    1972, 
    914.092975255705, 
    2277.79654107849, 
    2891.14299085074, 
    1368.01760643655, 
    1462.30419571459, 
    1442.55366504042, 
    2007.6770975194, 
    3168, 
    1994.00304396645, 
    2999.70286948908, 
    2150.12117886465, 
    2753, 
    1171.91441718416, 
    2215, 
    2374.58487809284, 
    2964.44576445461, 
    2021.90419562155, 
    2465, 
    1736.87740381559, 
    3084.82388991341, 
    2991.33750931652, 
    1409.45082545417, 
    1671.7149130801, 
    2466.54816540415, 
    1809, 
    2089.63073448677, 
    1578.87801849159, 
    1124.12694418139, 
    2896, 
    769.836581776866, 
    2390.53425127175, 
    1729.66103832228, 
    953.27384837633, 
    2611.78097901989, 
    2090, 
    2020.55106053113, 
    1784, 
    1335.30340757232, 
    2943, 
    2705.55422766163, 
    2077.05336603662, 
    2643.99852464651, 
    1345.88696599676, 
    2054.47642127526, 
    1308.31589187547, 
    2477, 
    2067.14206026275, 
    1784.22148954931, 
    2220.91216430245, 
    3070.73406703483, 
    1385.64225753029, 
    1319.60644231549, 
    1099.49676618215, 
    3113.04143788558, 
    1030.26930212565, 
    2744.07879121158, 
    1660.8836815165, 
    1950.50731553456, 
    2590, 
    1715.22259018577, 
    1011.59047657941, 
    1894, 
    635.644732629093, 
    2848.06447685511, 
    1152.94218486216, 
    3090.23898246713, 
    2573, 
    734.500794587833, 
    1943.12766145918, 
    2117.9001865245, 
    2311.74796051268, 
    2052.09360158491, 
    2431.3604700816, 
    291.721910558428, 
    1724.83249263333, 
    1179.00675603289, 
    1215.20751194372, 
    1674.42963813995, 
    2213.79529171975, 
    2819.49803502852, 
    1828.22386420334, 
    2141.88697681376, 
    1383.15259199664, 
    2628, 
    3132, 
    1565.56060381804, 
    1262.51566925237, 
    2489, 
    2554.81113903494, 
    1655.61315872205, 
    1969.01795175939, 
    2409.63393884343, 
    2433.99212479536, 
    958.601296420022, 
    1973.84098133506, 
    1776.22022990978, 
    875.793603104607, 
    1453.84046246451, 
    1886.92872003694, 
    2181.87899551045, 
    2838, 
    1767.49247453777, 
    2912.84198171106, 
    1379.45385473555, 
    2721, 
    2629.17634677199, 
    2709.84660497108, 
    1383.73810801472, 
    2158, 
    1296.79694794672, 
    1858.02978379001, 
    2893.75709750041, 
    2117, 
    837.07289632244, 
    2968, 
    3194.28921712437, 
    39.7213449022315, 
    2048, 
    3136.46383063669, 
    1290.71933496854, 
    2740, 
    2737.00695125313, 
    1624.22101558313, 
    1849.04043954148, 
    1913.19935343774, 
    977.091375400774, 
    2993, 
    708.940955195474, 
    2179.72019166845, 
    308.497486681239, 
    2071.74587153467, 
    616.043969126238, 
    1403.10714218498, 
    2819, 
    2956, 
    1079.52574967444, 
    1992.6536514013, 
    2722.07375361034, 
    2651, 
    1266.78422862359, 
    2277.57884104311, 
    1664.65913414327, 
    1367.89446172966, 
    2072.35744122392, 
    1146.87019572265, 
    2518.78532238603, 
    1780.2239211587, 
    965.271849073507, 
    2400.94269951058, 
    2882.74714680182, 
    2667.65574821054, 
    2149.38854123308, 
    3146, 
    58.4319936094383, 
    1845.21276307792, 
    1682.01352570063, 
    1755.78375153308, 
    1332.03392076409, 
    2904.53573978824, 
    1535.96438225634, 
    1019.07387185478, 
    856.161525751841, 
    2544, 
    1038.12478967938, 
    2663, 
    3163.91546095942, 
    1872.58572378274, 
    2105.7673134704, 
    685.805580332329, 
    2730, 
    592.348044581225, 
    1965.45259490399, 
    2264.41420248728, 
    376.396283012925, 
    1168.9996035627, 
    1500.83257842879, 
    2231.23244574699, 
    2747.01900218529, 
    1302.04843691969, 
    1847.34510273619, 
    2952.02645217953, 
    732.836235404459, 
    1885.61416026803, 
    2015.89106057055, 
    1227.8942367692, 
    376.172283718123, 
    2655.55893033931, 
    1765.19453548713, 
    1014.09240776995, 
    1058.66330022341, 
    1879.85150282889, 
    1900.81965501134, 
    3245, 
    1942.45344991771, 
    1775.55883730342, 
    1250.36815932935, 
    2958, 
    2070.83065623328, 
    2450.12710916266, 
    2778, 
    2009.51707368965, 
    1373.04185896731, 
    2526.33682500978, 
    2259.84609351649, 
    1659.09678316254, 
    843.252984643991, 
    2160.13016041223, 
    1578.01784861731, 
    3252, 
    1059.33101271091, 
    739.590598580477, 
    1145.17410985606, 
    1360.86552758274, 
    1970.48917050818, 
    1684.92173620243, 
    2623, 
    1349.64832372909, 
    962.440294894156, 
    937.679466374813, 
    2737.89690318297, 
    1868.27840906539, 
    313.714664913036, 
    2523, 
    1424.40698397745, 
    2446.45700532129, 
    2272, 
    2583.96945278868, 
    2756.91991257488, 
    2094, 
    2343.93463618885, 
    1316.0626097704, 
    1090.08013283759, 
    2105, 
    678.527594809112, 
    678.098808491651, 
    2337.00855313476, 
    3148, 
    2405.22352611094, 
    1134.25063134941, 
    2802.81574528162, 
    2948, 
    2513.14955922585, 
    1560.11460302216, 
    2003.20271478903, 
    2590.42164355054, 
    543.74177277436, 
    631.35734648173, 
    666.294043628362, 
    1587.13838664661, 
    3234, 
    2236.74168541969, 
    2312.78367016718, 
    2279.85183646626, 
    2077.26671094074, 
    1933.182031846, 
    1847.33103802442, 
    2764.02125688688, 
    2381.54232638654, 
    2351.23970220081, 
    1836.49047206241, 
    2960.09974656389, 
    3069.91709477401, 
    2764.423157993, 
    1874.37119934491, 
    1149.33171106362, 
    2751, 
    3035, 
    1955.36769146962, 
    1806.53704139065, 
    2027.60077921334, 
    2268.58106027656, 
    2008.09803526183, 
    2753, 
    2459, 
    2215.64428154866, 
    1587.13694610468, 
    1252.57661456266, 
    2520.5881942041, 
    2404.85523875012, 
    2587.5925972219, 
    2495.05744658287, 
    1987, 
    2496.40590962686, 
    2259.06367399268, 
    2906.80376919308, 
    1280.82699148558, 
    2644.33326790622, 
    1281.40046246164, 
    2546, 
    1210.838048117, 
    1555.59503631247, 
    1574.33895611673, 
    839.006157485803, 
    2025, 
    2161.75721515424, 
    3006, 
    3046, 
    2398.64823286246, 
    3199.60619417381, 
    1779.38849242511, 
    2533, 
    2461.51467555038, 
    2560.02962011684, 
    1429.14291149268, 
    2483.89418868039, 
    2184.25408350924, 
    2732.57361226037, 
    1383.00917561745, 
    1641, 
    1108.76689535621, 
    2225.87259103634, 
    1348.11929204594, 
    303.834939951865, 
    2868, 
    3114, 
    1558.23191222975, 
    2249.63165459227, 
    1464.79555288069, 
    1170.30948607616, 
    1916.80852344892, 
    1942.6999082431, 
    1807.08499873473, 
    1430.80361439287, 
    2920, 
    1731.42157635645, 
    1631.55699937243, 
    2636.34634787639, 
    2257.91059579551, 
    1383.80087498085, 
    1444.59416076574, 
    3000.0204501327, 
    568.507004782472, 
    1442.4743274576, 
    1128.64118021778, 
    1791.14760721962, 
    3080, 
    2837.98557276719, 
    1875.62850213326, 
    1859.8784927138, 
    2691.03362144731, 
    1965.74014101729, 
    2455.02813574548, 
    3124.73701174329, 
    1195.97562264213, 
    2523.40217324055, 
    1900.35947184005, 
    2941.63792871637, 
    2546.62691528062, 
    1153.95414710749, 
    2270.50228484001, 
    2073, 
    2451.05334043658, 
    1259.74140166099, 
    1154.88328576468, 
    2982.90919292801, 
    716.46301005515, 
    1054.4365478169, 
    838.674442832968, 
    1197.62516776942, 
    2112.39207054911, 
    1201.60311672756, 
    2231.54596029549, 
    1852.99013656459, 
    2385.61099306815, 
    1800, 
    1763.48499706052, 
    1976, 
    1938.56141905756, 
    3075.32279399592, 
    1999.35258111801, 
    2781, 
    1643.95279780012, 
    2370.5649756195, 
    2559.79984473891, 
    2259.35270251036, 
    2061.07685599653, 
    1653.79997975232, 
    1207.64122363233, 
    3195, 
    1001.81056619515, 
    2857.45637889117, 
    1888.95525489165, 
    1355.62175648186, 
    1555.09802057433, 
    2274.25491848208, 
    2009, 
    1292.96064295414, 
    2251.30034116468, 
    1910.30860045329, 
    972.037279972797, 
    2978.08802605834, 
    2531.96983186056, 
    1345.53382912207, 
    1531.66812487372, 
    966.218724342211, 
    2193.62903985839, 
    1991.00370730543, 
    2156.09833165964, 
    2155.01882590309, 
    1112.12012787201, 
    1730.7607067935, 
    1995.11174369796, 
    1320.16975973459, 
    2114.69887159107, 
    1633.05585076189, 
    2532.72180453888, 
    3142, 
    680.312612479362, 
    2690.80014406818, 
    2728.40274274922, 
    1287.7018136261, 
    2214.67529744329, 
    2184.7998067837, 
    1306.23673384486, 
    2243.39748958148, 
    1384.18998926215, 
    2057.99041308686, 
    2762.47594500096, 
    1625.27996847405, 
    3073, 
    1476.3019421666, 
    1111.03089406047, 
    2582, 
    2571.18221684131, 
    2521.04801339414, 
    1586.0511248394, 
    1802.94764238701, 
    1754, 
    2605.51527133467, 
    1108.68362846577, 
    2777.61395626991, 
    1608.34336621792, 
    2115.95420020187, 
    1430.12560140134, 
    2486.66132075333, 
    2977, 
    3227.94154243763, 
    916.681118394941, 
    3010.65100002615, 
    2808, 
    2874.49047667836, 
    2273.27776824072, 
    1641.24609300187, 
    1000.63284861753, 
    2049.78010808242, 
    1385.6023435034, 
    1363.66235504459, 
    2949, 
    1421.67511309036, 
    2376.55193865069, 
    1340.78338404406, 
    1815.24274383907, 
    1226.13886171471, 
    2342.18736584984, 
    2701.64290090851, 
    2842.33269150185, 
    2033, 
    2563, 
    3033.99465419402, 
    1321.08354423552, 
    1433.79310349048, 
    2470.54397647722, 
    1654.23236425969, 
    1041.19553248807, 
    2046, 
    1416.33155085196, 
    1874.28913543732, 
    2693, 
    2976, 
    2832.07361993487, 
    881.351265343466, 
    2437.35569920353, 
    3201.06245489827, 
    2181.18971064732, 
    2061.24115947479, 
    2781.29515704762, 
    865.150902577699, 
    2118.46073356335, 
    1358.56755742795, 
    847.994961421305, 
    2440, 
    1132.65327643864, 
    1635, 
    2757.2101943427, 
    3165.90170373171, 
    1553.48546684702, 
    1779.78213836517, 
    2129.28791492061, 
    1050.13887518712, 
    2034.66135187898, 
    1189.84091288141, 
    2132.96508197937, 
    1955.82323630545, 
    1607.1987902662, 
    2945.1090077821, 
    1813.52124767538, 
    1881.52723506061, 
    2319.93478059634, 
    1716.10717314963, 
    2422.78679058906, 
    2800, 
    1253.81340329283, 
    1627.96263983182, 
    1628.94995960228, 
    2028.96978604992, 
    3215, 
    108.797730587061, 
    3022, 
    2137, 
    771.193532984451, 
    2783.0048015092, 
    2536.71001491443, 
    43.4171948535668, 
    2352, 
    2335.2893675356, 
    2498.63277032051, 
    1607.64418651441, 
    2366.97390982076, 
    1584.39269302331, 
    3160.15737885204, 
    1175.17071353899, 
    3050, 
    2372.02578766947, 
    1911.87773664908, 
    2574, 
    1600.14621790744, 
    1771.21000855146, 
    1741.53949370688, 
    869.301182118135, 
    2801.64635550486, 
    733.306160366054, 
    876.568816342765, 
    2547.02276556707, 
    802.682316297247, 
    1973.36440740352, 
    2662.26225179458, 
    1029.6629445037, 
    2243.62599665026, 
    2154.60185225237, 
    1425.29235886182, 
    2846, 
    2825, 
    2085, 
    2530.49272919579, 
    2355.2072550528, 
    879.883791794999, 
    2260.57500657718, 
    3117.99754319773, 
    1863.85319294434, 
    1260.83727692768, 
    2324.3705395212, 
    3048, 
    919.433307067185, 
    2656.52334725904, 
    2745.47860617025, 
    1404.3104023921, 
    2854.58349488262, 
    3158, 
    2471.33763376701, 
    2115.99007114513, 
    2047.92534311478, 
    1447.67511492592, 
    2080.4309422335, 
    1980.35854207215, 
    2574.92263063053, 
    816.626348766627, 
    2006.91862474966, 
    1460.36797619052, 
    1211.30052457752, 
    2787.03678246038, 
    2935.80049963329, 
    2538.05684617156, 
    2684, 
    3104, 
    2058.2252622813, 
    1023.0720913185, 
    2398.08339346107, 
    1720.67087425278, 
    2578.96360111195, 
    2199.18747016149, 
    2088.81830992242, 
    1630.36838325195, 
    1602.70197275168, 
    2999.23344911815, 
    2133.38264042286, 
    2355.56038921137, 
    2699.04529376075, 
    1849.91032879368, 
    2769.82374080505, 
    1803.06662998425, 
    2805.79144109992, 
    2179.80574077902, 
    2816, 
    1235.54923522901, 
    2353.48128251713, 
    1015.39330779461, 
    1001.62096123151, 
    2667.64431320493, 
    1922.82982355403, 
    2100, 
    1739.32980303409, 
    2976, 
    3142.03400989879, 
    2200, 
    3177.75893890449, 
    2677.96147443844, 
    2644.27376193478, 
    3008.23666420169, 
    1401.13411242463, 
    2207.02215274222, 
    1264.34294547046, 
    2924, 
    1493.35347953119, 
    2000.76444474547, 
    2150.68021376291, 
    693.785803629985, 
    2865, 
    3028, 
    1301.44605390785, 
    1701.57599602744, 
    2467.80031213461, 
    2543.01897080417, 
    2891.81447717316, 
    2145.74281442774, 
    1778.94334708672, 
    1983.64008771931, 
    2819, 
    1718.3925230007, 
    2107.13728123665, 
    2799, 
    2531.35767449504, 
    1297.9896473722, 
    1925.59975805898, 
    3091, 
    1192.33972021742, 
    1488.29863809933, 
    1391.76605039795, 
    1886.50373757044, 
    2980.81608203869, 
    2772, 
    2592.78904883883, 
    1670, 
    1412.84960791786, 
    2602, 
    1143.49030178708, 
    1533.63990790725, 
    2591, 
    3158.11966378168, 
    1177.32685144962, 
    2328.80640082772, 
    1352.40897877209, 
    2865.09011511004, 
    756.618452783949, 
    1467.61194562165, 
    1394.58916389581, 
    1924.0000421797, 
    2217.62493528049, 
    1736.929585882, 
    2984, 
    1753.47427434952, 
    2488.68490328571, 
    1446.36415206534, 
    1323.25328114558, 
    1995.25134582401, 
    1666.17001900639, 
    3189.21518970848, 
    1880.89085427123, 
    1339.59869151315, 
    2895, 
    1951.01174243567, 
    1079.1692005325, 
    1603.58875680831, 
    2489.7334804894, 
    918.793378984655, 
    2001.27855436596, 
    1586.05551140307, 
    3261.52091769947, 
    1047.446896814, 
    2951.80913054529, 
    1921.09292832432, 
    1742.97078168259, 
    63.0745204287434, 
    1854.43407710944, 
    2047.45489073255, 
    1616.59715176943, 
    2504.08642721212, 
    1077.84669878765, 
    2840.36473593633, 
    1016.0014235222, 
    2418, 
    1713.7537165135, 
    2549, 
    2245.40435754819, 
    1584.8624881108, 
    1126.98003976153, 
    2468.80225335439, 
    2017.15554321202, 
    2199, 
    2393.17473416214, 
    3140, 
    2095.54352068057, 
    1284.9970884882, 
    2855.4306213108, 
    2865, 
    2404, 
    2463.58750780051, 
    1899, 
    1245.59266503061, 
    530.896922534884, 
    1392.2068128703, 
    1520.526710879, 
    1479.30914272348, 
    3184, 
    1946.04562533048, 
    2427, 
    2435.63743027206, 
    2320.13682918195, 
    1789.81844797801, 
    1823.94889904768, 
    308.316258986418, 
    2620, 
    2165.9708473362, 
    2994.32813103491, 
    3149, 
    2787, 
    2971.97400210363, 
    2360.21822256809, 
    2416.83201742767, 
    1767.71964467615, 
    2846.79306026279, 
    2525, 
    2039.05787440838, 
    1296.10751992596, 
    1167.86546620243, 
    2080.37702105509, 
    2540.03671660115, 
    2704.68864113653, 
    2303.53195854623, 
    2033, 
    2108.43277363291, 
    2398.49237101447, 
    1527.85708938825, 
    2964, 
    2406.94999506582, 
    2604, 
    1519.8110465947, 
    1827.92864122245, 
    1134.69142469381, 
    1962.21366112074, 
    2658.77488573607, 
    3015, 
    2968.18608142911, 
    2509, 
    3203.05884844985, 
    797.741947465438, 
    2430.02129764915, 
    2324, 
    1973.37064232008, 
    1707.6032242524, 
    2620.76019494725, 
    1079.57301715392, 
    2735.19301578955, 
    1886, 
    2375.0353324965, 
    1445.17167096524, 
    2310.52401221985, 
    1396.9220064516, 
    643.959636669324, 
    2832, 
    3155, 
    2315.58507020239, 
    1696.43492043352, 
    1678.56966824598, 
    2025.33259116804, 
    2053.83737719239, 
    1673.10773886762, 
    1340.93412960598, 
    2920, 
    1665, 
    2526, 
    2926, 
    722.640410690814, 
    1524.47363095108, 
    1333.63882247029, 
    3142, 
    2956.64639662802, 
    1992.82454709579, 
    2061.65981054315, 
    2732, 
    2133.63729077497, 
    2410.66863493382, 
    2510.41417286195, 
    1777.90146432009, 
    3038.91258320731, 
    2947.5667517389, 
    2530, 
    2401.60217961417, 
    1880.57904815889, 
    2933, 
    1694.04756378849, 
    1927.99611495675, 
    2000.83677038122, 
    1894.93182118366, 
    2994.46403027597, 
    2638.74214181908, 
    2067, 
    1322.53452054172, 
    2687.78424681025, 
    1449.69130672255, 
    1917.76299591929, 
    1953.18990043485, 
    3013, 
    1443.21086818591, 
    757.491869360356, 
    3137.93476749307, 
    1072.30605715246, 
    2786.34743476289, 
    1524.04982920048, 
    1298.58728277549, 
    1086.08430663935, 
    1058.4649718575, 
    2804, 
    3057.25345138496, 
    2606.64209757639, 
    1825.76969602516, 
    1839.09518548607, 
    2095.93547339157, 
    2379, 
    2090.02956629595, 
    2352.57939885067, 
    939.896918901097, 
    1798.26648913993, 
    1786.54152187466, 
    2781.48776895095, 
    1624.38524585116, 
    401.459457566284, 
    2185.98924353941, 
    1376.1852686997, 
    2599, 
    3140, 
    1122.65178059417, 
    2552, 
    2034.79691092592, 
    2063.59043567006, 
    2363.32044467149, 
    1718.80684816694, 
    1208.00330575016, 
    3055.63665417086, 
    1755.82012036524, 
    2046.23953354466, 
    2874.48027792277, 
    1727.06822678867, 
    2972, 
    2673.62203442189, 
    2647.28423293968, 
    2661.4632600149, 
    1440.74989267382, 
    2083.40257697416, 
    1486.14007806891, 
    2030.45256086374, 
    2420.51716504905, 
    2962, 
    3220, 
    1952.05322501151, 
    3111, 
    2767, 
    2786.5014597282, 
    2483.58591422133, 
    1636.37760483449, 
    1626, 
    738.900101136043, 
    2989, 
    2259.80154507805, 
    2063.28886800595, 
    2780.95796473967, 
    2925, 
    2039, 
    1146.27693939114, 
    3023.92899904077, 
    2342.07054393057, 
    1623.0170367151, 
    2079, 
    2012.60521645019, 
    1818, 
    1330.83754424094, 
    2526.98078944336, 
    2918.74526171279, 
    2725.80476784136, 
    2275.76733352566, 
    3169, 
    513.383675052567, 
    1990.08112085959, 
    1853.33175993542, 
    1024.51070025649, 
    2870, 
    815.719667670785, 
    2041.51202226141, 
    1750.20175942693, 
    2511, 
    2705, 
    3166, 
    2615.90687838834, 
    2187.5760922396, 
    1213.02754245613, 
    1216.46569476674, 
    2203.03124452032, 
    1870.82463330647, 
    2950.49402237511, 
    1117.24666928942, 
    2130.23673458327, 
    2705.23042832474, 
    1527.40873589943, 
    1169.75904657547, 
    1799.88431629774, 
    3255, 
    1752.7603950081, 
    2985.52402289047, 
    975.298708940675, 
    2793.05569596232, 
    2331.6023978819, 
    2471.34660125219, 
    2268, 
    1884.38775004726, 
    2242.87432506032, 
    1530.91658085447, 
    3232, 
    1093.29500221573, 
    3024, 
    2218.06057569767, 
    1097.54788221368, 
    1193.34231792908, 
    1901.81854573007, 
    2688, 
    1030.06700776759, 
    993.05649448979, 
    2677.56353659292, 
    629.961191357346, 
    1298.88686111342, 
    2384.78456485848, 
    2244, 
    816.745235030274, 
    2654, 
    2838.04443354244, 
    2404.49931377995, 
    1113.42600330772, 
    2328.23785057219, 
    3147, 
    2006.97593997704, 
    1164.92306882979, 
    2686.54021446018, 
    2983, 
    2559.384812287, 
    1382.59645826448, 
    1239.49911830274, 
    2532.19985855873, 
    1531.44524434987, 
    3214, 
    2330.94932277479, 
    2247.49223782199, 
    2224.22928493628, 
    1876.86984753712, 
    1880.68572690082, 
    2708, 
    748.290146290137, 
    2270.12265814065, 
    2928.5152808703, 
    3026.51221661453, 
    2699.56872717548, 
    2736, 
    3061, 
    2072.65028280199, 
    1479.94700390994, 
    2102, 
    2704.31111750781, 
    704.135374962166, 
    2375.43022157389, 
    2259.49920159176, 
    2319.69770597437, 
    2510.0445744045, 
    2565.35571512658, 
    1944, 
    2605.05350122146, 
    2148.3869125084, 
    2880, 
    2489.76035303904, 
    2054.85417418094, 
    2991, 
    3081, 
    2336.86980059125, 
    3193.59743319981, 
    2583.3854083723, 
    2544.96939082686, 
    1201.66044861344, 
    2827.03766744374, 
    1766.56648141821, 
    2190.97878948771, 
    2881.70662345429, 
    3089, 
    1142.35415400725, 
    2743.73813040854, 
    789.934290307124, 
    1830.31019478583, 
    1954.08107253409, 
    1889.21698978933, 
    1865.62116644124, 
    2890.2262012761, 
    1684.02273014543, 
    2694.02220428108, 
    2376.09520919549, 
    1416.79556387646, 
    3035, 
    1051.45814058746, 
    3051.85651448215, 
    1747.13570189374, 
    583.379881296564, 
    2663, 
    1856.02955454434, 
    2499, 
    2469, 
    1866.6570681751, 
    2923, 
    2502, 
    2150.19702221821, 
    2126.28145113034, 
    2997, 
    1219.40988272321, 
    1042.66364357683, 
    2332.56990438087, 
    1700, 
    1984.68565484512, 
    1707.24024718012, 
    3121, 
    2429.33285188548, 
    1962.25743629916, 
    2821, 
    1769.51277289715, 
    2468.42487468518, 
    1226.59635923576, 
    1796.78262074414, 
    1388.35921737914, 
    3218.15969437892, 
    983.478759386983, 
    2891, 
    1396.46851374014, 
    2936.36631534407, 
    2456, 
    1347.92888613091, 
    2283.61600274828, 
    1924.62364989441, 
    2553.42974141286, 
    2187.9020616978, 
    1971.3450720616, 
    1850.28296446063, 
    2074.9194314754, 
    2389.21203103114, 
    1771.44225629301, 
    2494.94844918968, 
    3141, 
    2748.91314339457, 
    2777, 
    1755.40641947624, 
    2273.22607339674, 
    2088.4204692495, 
    1808.67130134377, 
    1166.02690957849, 
    2627.43052837774, 
    1524.7708807627, 
    3114, 
    1621.93395925365, 
    2532.33354063212, 
    2533.08624719519, 
    2457.8674051326, 
    1805.3484493266, 
    1076.10445739944, 
    2741.79860026431, 
    1493.50219379139, 
    2985, 
    3207, 
    2807, 
    2910, 
    1362.16960198016, 
    2597.33488258269, 
    1951.38800168497, 
    1503.30301975774, 
    2921.90157278117, 
    2444.77562922642, 
    1857.07057932016, 
    1881.81663603657, 
    1324.87976787022, 
    2654, 
    2797.7846704046, 
    2019.8484134217, 
    665.486357286462, 
    1414.33366080395, 
    2519, 
    1646.99216728936, 
    1126.74303820887, 
    115.755573353661, 
    1904.54761032313, 
    3000, 
    2880, 
    3204.03312298946, 
    2155.8638753283, 
    1558.1099378034, 
    2400.14283949682, 
    1225.19043216463, 
    2786, 
    3164, 
    1735.66892109081, 
    1939, 
    1367.37754979618, 
    2095.50522389877, 
    2931, 
    1741.84132833808, 
    2847, 
    1321.62941121172, 
    3194, 
    3024, 
    2768.62743245781, 
    2288.11414284952, 
    2360.4371146308, 
    1640.38578464098, 
    2416, 
    1672.0134612191, 
    3132, 
    2525, 
    1960.73694069563, 
    2850.72030595228, 
    836.299724160816, 
    2481.29156894036, 
    769.825754679287, 
    2175, 
    1653.31331221879, 
    1220.72184965211, 
    2898.85472047732, 
    2772, 
    2582.5388676003, 
    1168.83576847003, 
    2481.63404814349, 
    800.234169401291, 
    2245, 
    1238.90893157561, 
    1955.07060036041, 
    3077, 
    949.982779729653, 
    2700.96432187059, 
    1935.7984525468, 
    972.200874345116, 
    2899.64114269882, 
    3128, 
    2525.85743759326, 
    2015.11773432455, 
    2019.27218217355, 
    2508.5467587988, 
    1895.41275200926, 
    1433.25828044403, 
    2629.280086305, 
    2883.29753819627, 
    2331.30610592076, 
    801.967971914674, 
    2651, 
    3117, 
    1670.53240982929, 
    1841.44895916315, 
    2340.13319994149, 
    2510.24299272043, 
    2104.35654762528, 
    2037.75538345354, 
    720.77472421114, 
    2035.2251076471, 
    2272.69495347947, 
    2764, 
    1802.42426411586, 
    2848.3511147862, 
    1650.09066845607, 
    2764.15625531785, 
    2403.75676438275, 
    2778.19840121592, 
    2266.08734109528, 
    994.870000358102, 
    2290.96069888594, 
    2978, 
    3170, 
    3165, 
    2699.51244277807, 
    2966, 
    2093.97289404207, 
    2108, 
    1134.67922459658, 
    2847, 
    2999.89840875289, 
    1891.11434913182, 
    2428.76281825759, 
    2210.31717905764, 
    1724.53720419426, 
    2035, 
    2723.97967376441, 
    1739.64636641332, 
    583.626942776793, 
    2842, 
    2598.50671049267, 
    1173.54207916749, 
    3122, 
    1636.05769877153, 
    2948, 
    1270.16176190566, 
    611.385832847031, 
    2571.7657350903, 
    1785.39216295947, 
    2635.61917322734, 
    3160, 
    1142.88217445012, 
    2779.68118476806, 
    829.262626983324, 
    1230.46053103808, 
    1071.19192788403, 
    1759.67120120235, 
    2242, 
    2972, 
    1573.14786312592, 
    333.330598581993, 
    2577.97234568006, 
    1290.22829889507, 
    1951.7147766698, 
    1796.31731640404, 
    3225.29623215394, 
    1839.89984519813, 
    1272.36043791504, 
    2930.99506703353, 
    2516.38313049338, 
    2545, 
    2181.45969413263, 
    2085.5248271064, 
    1611.32581597722, 
    3273, 
    1048.05049532861, 
    75.5932052844959, 
    2025, 
    1715.52543503925, 
    2566.43839152718, 
    1041.67443675978, 
    2793.67034121963, 
    1586.34905318109, 
    2501, 
    2266.03783803249, 
    2099.69561663611, 
    2651.69131739921, 
    2282.80223644703, 
    1051.32440127798, 
    1265.62995009216, 
    1195.20620707852, 
    2380, 
    3140.35998991344, 
    2866.6925710289, 
    2902.85821753034, 
    353.992012933982, 
    2463.18268593662, 
    1768.40306629375, 
    1877.83137980056, 
    2366.0138816775, 
    528.177345199646, 
    1677.15697241123, 
    1580.72239236874, 
    3211.27274304122, 
    2104, 
    2365.71487414995, 
    2392.74465791935, 
    2224.67842357039, 
    1832.92376307156, 
    2821.5613974576, 
    2997.84632159301, 
    3113, 
    2769, 
    3005.46851057873, 
    2363.30357649715, 
    1900.63012915158, 
    2799.02535016182, 
    2515.0593314888, 
    2183.09449676862, 
    1472.14285963875, 
    1062.24664163569, 
    2478, 
    2652.12208830394, 
    2413.23376647714, 
    2018, 
    2350.32892288433, 
    2324.63723450692, 
    2939, 
    2587, 
    1400.5441471213, 
    1986.99227544965, 
    2481.32491107383, 
    3011.92241657576, 
    3004, 
    3196, 
    2400.05997492051, 
    2353.07306052234, 
    1744.09769792302, 
    2589.51563979864, 
    1549.83590052416, 
    1550.53119556851, 
    2276, 
    1441.66284808585, 
    440.36832043864, 
    2851.93260333092, 
    3137, 
    531.505725675977, 
    1570.98475418857, 
    1450.84584860714, 
    485.137394945705, 
    1982.47612382674, 
    1732.5744452806, 
    1475.69583029002, 
    2915.89146307684, 
    1747.20018910349, 
    2579, 
    2208, 
    1255.88649868391, 
    2961, 
    986.016847916532, 
    674.251639743187, 
    3112.2321780801, 
    1084.00370708959, 
    2911.99440130208, 
    1965.1673390638, 
    2713.877553587, 
    2058, 
    2455, 
    2554, 
    1863.27831532873, 
    3000, 
    1335.77267602593, 
    2570.33431239374, 
    2199.56985317369, 
    2330, 
    2337.56083085558, 
    2957, 
    1693.78078062109, 
    2104.04400312717, 
    1685.11914943172, 
    1910.45766910827, 
    1959.02771551528, 
    3036.97905421681, 
    2034.05280069731, 
    2735.10457181909, 
    1543.2803573918, 
    2015.34149908777, 
    1546.8612783598, 
    3167.8417848924, 
    1058.00599533206, 
    2826.75520034206, 
    1189.77899102628, 
    1458.86532188122, 
    958.552492858217, 
    3017.86478784685, 
    2573, 
    1691.51295520703, 
    2044.73501079985, 
    2122.10273385262, 
    2274, 
    1923.65917514273, 
    2568.55778474824, 
    3141, 
    752.506602162741, 
    2621.68983184633, 
    2132.12452148983, 
    2272.57972694875, 
    1428.19847117311, 
    986.253562071756, 
    1516.25758222055, 
    1877.967829681, 
    2860.6857569676, 
    1676, 
    3031, 
    2627.37088285724, 
    2597.96170780731, 
    2593.11186894573, 
    1939.31836170949, 
    1650.27159505745, 
    1474.48495160124, 
    2968.33890450083, 
    3234, 
    3069.96295996637, 
    832.474980437224, 
    2793.02741036892, 
    2831, 
    1642.37815421343, 
    1100.50285195618, 
    2976, 
    2323.13869356645, 
    1997.14865223587, 
    2740, 
    2887, 
    1731.56693962855, 
    2036, 
    1618.00353124057, 
    2073.09167618533, 
    1863.38219043875, 
    1839.61450291211, 
    2950, 
    2779.80294419106, 
    3187, 
    1923.15603823354, 
    1710.53544023254, 
    2824.37535072108, 
    2119.32962302597, 
    2519.13046540204, 
    889.343908664669, 
    970.43367275368, 
    2474.98889920142, 
    2733, 
    3166.9337442074, 
    1800.67657555858, 
    2417.17916554817, 
    2116.9040055332, 
    2166.62897674471, 
    2940.79426545821, 
    1659.64039763988, 
    2754, 
    1456, 
    1251.56110006223, 
    1794.01022013539, 
    3237, 
    3009, 
    2794, 
    1829.02558216552, 
    2417.25887889922, 
    2288, 
    2136.0244463212, 
    2301.40626556525, 
    1529.22091797244, 
    3201.31988162449, 
    1115, 
    1254.02547652788, 
    1360.23362123104, 
    1524.41920356775, 
    2745, 
    2522.50198693757, 
    2654.64284472424, 
    2631.97934130178, 
    3197, 
    2627, 
    3112.88322996232, 
    2129.19340341477, 
    2576, 
    2651.04111421673, 
    2724.68304018013, 
    3006, 
    1839.65721510533, 
    2697.92238621414, 
    2347.67646271063, 
    2917, 
    2492.94730795613, 
    1667.96859411156, 
    2489.06892857468, 
    1124.98161796861, 
    2754.51754021202, 
    2435, 
    2472.57519699772, 
    2008.67782129179, 
    2771.33629188393, 
    3145, 
    2469, 
    2382.92653038912, 
    2762, 
    2773, 
    2708.77587602071, 
    1895.61636857079, 
    614.379198759562, 
    2754, 
    1848.49142892978, 
    1087.04884374572, 
    2372.54118715055, 
    2224.30015547961, 
    1645.90283281041, 
    2554.61055924517, 
    2494.16544015411, 
    2884.23624213479, 
    1977, 
    2302.7876999352, 
    3171, 
    2604.0963121064, 
    2872, 
    1798.33251832983, 
    2444.80780557747, 
    2642.99803248502, 
    3061, 
    814.584615682059, 
    3175, 
    2640.1940316125, 
    2672, 
    3093.11393971183, 
    1220.43506773575, 
    1808.35952919302, 
    1319.46149798863, 
    2133.22919691364, 
    1186.43282486429, 
    1918, 
    2095, 
    2110, 
    1831.58898902809, 
    1788.539676332, 
    2896, 
    2574, 
    2547.6670477385, 
    1495.43382744517, 
    1784.17852579724, 
    1903, 
    2179.59231583636, 
    2781, 
    3020, 
    3027, 
    1541.2091783847, 
    2826, 
    2097, 
    2617, 
    3036, 
    2058.5226089672, 
    2569, 
    2980.91087856332, 
    3056, 
    2522.71681066029, 
    3061, 
    1872.16850432681, 
    979.40264330763, 
    1961.82788876687, 
    1760.54708944243, 
    2863, 
    2294, 
    2632, 
    1843.65417276635, 
    1760.25485703311, 
    3041.22854464078, 
    2228.54604377039, 
    2774.79523342792, 
    2882, 
    2289.98818549024, 
    2682.7566094322, 
    2140.58399499815, 
    2264.21037595965, 
    2495, 
    2223.51456826734, 
    1892.07551160952, 
    2717, 
    2457.95073029208, 
    2514, 
    2962.72536791912, 
    2269.28701251433, 
    2384.88620592948, 
    1729.62049832335, 
    1895.39591234035, 
    2270.82938810093, 
    1983.74035784081, 
    1976.46077779498, 
    3189, 
    1216.1480906, 
    2383.89971513514, 
    1670.55819817851, 
    2616.25737855017, 
    1850.97813699242, 
    3086.44813459961, 
    3278, 
    1654, 
    2797.17703227592, 
    2457, 
    3120.31743249524, 
    1964.14883127815, 
    2970.14139057441, 
    2862.15031255082, 
    2458.66636082748, 
    2643.36704117033, 
    1906.21258291158, 
    2155.53393244323, 
    1692.15043474167, 
    2938.98716713111, 
    2159.04590936773, 
    2835, 
    2926.32008837125, 
    2811.99848574678, 
    2605.14511200852, 
    2261, 
    2940.37438099506, 
    2158.0669167223, 
    3116, 
    2811.28441866499, 
    2148.62027827923, 
    3019, 
    2033, 
    2606, 
    2766.73907251886, 
    2861, 
    2203, 
    3154, 
    1508.78260129205, 
    2643.96178671663, 
    3049.64143661176, 
    2076.21052234087, 
    2556, 
    1546.48169519749, 
    2684.23477454345, 
    2526, 
    2813, 
    2937, 
    2622.81392471722, 
    3030.19587089412, 
    2170.92205242779, 
    2658.52062445814, 
    764.305568339152, 
    2279.46866808163, 
    2769.38272397372, 
    1535.01961130962, 
    1735, 
    2185.50160176819, 
    2226.95497422306, 
    1515.9246177712, 
    2723, 
    2967, 
    2156, 
    2382.10702671869, 
    1621.8168920027, 
    2754.32192117752, 
    2122.00323160389, 
    2459, 
    2382.41657624635, 
    2845, 
    2556.12736830835, 
    1921.38555628273, 
    2124.57317498856, 
    2421, 
    2455.28164791414, 
    2951.06535367057, 
    997.729929631794, 
    2873.03225071376, 
    1580.35710445194, 
    1116.86269673033, 
    1965.84655066229, 
    1966.83876808337, 
    1860.05698965512, 
    2852, 
    2836.95924147543, 
    1173.74889906494, 
    1200.66339651981, 
    3009.69989080351, 
    1399.58692293768, 
    1401.97238401049, 
    2290, 
    2782.74155062531, 
    2919, 
    2459.04638141891, 
    2069.73483098643, 
    3023, 
    1903.54783662203, 
    1754.65303661236, 
    3194.79060932354, 
    2990.45717024628, 
    1384.65961206062, 
    1966.79577221076, 
    2512.6252855432, 
    2690.64330331663, 
    2664.93369981231, 
    2450, 
    3164, 
    1848.75502008869, 
    3093, 
    1905, 
    1175.61526680351, 
    1919.77519560091, 
    933.522119998021, 
    2106.69835241879, 
    1598.77445640759, 
    1633.20854201165, 
    2491.98788965065, 
    2806.44546679182, 
    2872.28407637207, 
    2121.28911695822, 
    3185, 
    1451.02115389261, 
    2046.5278162903, 
    1896.41454818841, 
    2228, 
    3006, 
    3113.15233446514, 
    2648, 
    1206.77020262408, 
    1581.14412738903, 
    2415.54349156191, 
    2467.45228361111, 
    2951.97577576111, 
    1941.1232416891, 
    2582.91584712039, 
    2529, 
    1494.79999171173, 
    1711.91313229807, 
    2296.96918929667, 
    2858.42719012178, 
    2592.36437313641, 
    2278.81252833914, 
    1409.91947162014, 
    2141.95813627865, 
    1950.27512728866, 
    2512.9968554174, 
    2168.91949922319, 
    1931.60782263545, 
    2659, 
    2830, 
    2233, 
    2978.06532520491, 
    2644.33059954412, 
    2514.66731586441, 
    1675.65463267965, 
    992.612537380537, 
    2997, 
    1690.78555717787, 
    2234, 
    2546.82957849506, 
    3123, 
    2088.43041509187, 
    1828.83407003201, 
    2819.28318792913, 
    2949.80760126632, 
    2977.49147773657, 
    2533.68842884298, 
    2620, 
    2858, 
    2751, 
    1725.42441263875, 
    1876.88748989874, 
    2896.78928178098, 
    1683.62208541212, 
    1994.02502190338, 
    2511, 
    2668, 
    2310.747807218, 
    795.785735070254, 
    1816.15058526119, 
    1836, 
    620.054502371582, 
    1272.33076117416, 
    2141.67763640638, 
    2038, 
    2232.00081704792, 
    2488.47933722348, 
    2197.55924165553, 
    2848.25239961821, 
    2609.60793709837, 
    2499, 
    3232, 
    3193.90807137145, 
    2588, 
    1838.21468375436, 
    2871.72161768675, 
    811.286216900206, 
    2583.61721401187, 
    2262, 
    1911.03551375143, 
    3276, 
    2472.29628866514, 
    2453, 
    2287, 
    2251.56217114263, 
    2958.44474801276, 
    1561.56179298703, 
    2829, 
    2483, 
    2753.43021495267, 
    2369.2335355762, 
    1998.25843128391, 
    2200.09890074243, 
    2957, 
    2172, 
    2812.7624608466, 
    1478.53911551649, 
    1290.2421785013, 
    2636.37180507733, 
    2588.67700583008, 
    2268.38575533432, 
    2687.03820628296, 
    2757, 
    2620.51054818952, 
    1730, 
    3087.24472295127, 
    2486.19040333939, 
    2375.49355061268, 
    1900.14780070752, 
    2534, 
    2305, 
    2750, 
    2675.0661382623, 
    1368.88534523841, 
    2831.99521550085, 
    2311.08510150803, 
    1569.50253258159, 
    1213.46654167155, 
    2218, 
    3079, 
    2037.97109526576, 
    3013.02963227951, 
    2935, 
    2522.46894387112, 
    1390.86923294301, 
    1781.43477149195, 
    3107, 
    2123.67243676264, 
    2011.48147212578, 
    2169.78997436011, 
    977.853906588677, 
    1912.81728362995, 
    2977, 
    2353.70702688691, 
    2686.51493362753, 
    2582, 
    2844.904823745, 
    2782, 
    2819, 
    2904.01844708742, 
    2379.29112337841, 
    1713.01319102045, 
    1466.26221620583, 
    2776.34931270836, 
    2809.99390994874, 
    1834.88970280325, 
    2308.32572676156, 
    2204.24024936606, 
    2342.96578961266, 
    1783.98225709455, 
    1484.0913382417, 
    1734.65914378158, 
    2548.69646738227, 
    2385.88367798922, 
    2757.55059517135, 
    3231, 
    2826.63123789085, 
    2114, 
    2666.42279396959, 
    2269, 
    1844, 
    3092, 
    2153, 
    1528.95896885549, 
    3205, 
    1607.11731650097, 
    2563.524603888, 
    2542.02856464819, 
    2684.38270009874, 
    2484.50790856399, 
    3033.92205233005, 
    2847.1559764928, 
    1794.05372861604, 
    3128, 
    3142.04663824819, 
    2256.62960263857, 
    2511, 
    2892.97124462876, 
    3016, 
    2294.86048652823, 
    1502.02834121767, 
    2521.80029982752, 
    2476.3645474331, 
    2601.73634612163, 
    2490.38797933872, 
    2643.76733506579, 
    2570.36867259735, 
    3097, 
    2129, 
    1268.75136917914, 
    2568.99118054399, 
    2858, 
    1835.29088574854, 
    3006.62307657432, 
    2325.39473716912, 
    2540.53243814565, 
    1900.86271198698, 
    2469, 
    1302.40099421058, 
    2739.97830960954, 
    2403.31274410792, 
    2538, 
    1957.45118030926, 
    2829, 
    3165, 
    2059.3890007619, 
    2764, 
    2908.15920652238, 
    3103.81032348086, 
    866.732583679802, 
    1964.0115963527, 
    1161.74226099315, 
    2473.69631980845, 
    1222.07991913354, 
    2686.50618149488, 
    1659.10779526212, 
    2545.30343119413, 
    2496.11067800601, 
    2458.91236250901, 
    2884.54763347705, 
    2036, 
    3165, 
    2607.40051930308, 
    2845, 
    1792.69014009088, 
    2483, 
    2605.06881714796, 
    3067, 
    1237.72343866765, 
    3179, 
    2703.84648590492, 
    2644, 
    3073, 
    1710.63503206523, 
    1474.11601586182, 
    2113.89986866785, 
    1427.60184194491, 
    2107.11448475797, 
    2062.09704163383, 
    1738.82670606159, 
    1843.43357798955, 
    2871.79415595304, 
    2581, 
    2496.17390310169, 
    2572.33398046095, 
    2253.10068305699, 
    2783.06284381764, 
    3016.9032689658, 
    3045.65632924587, 
    1426.88032536099, 
    2853.09314754045, 
    2068.78941688456, 
    2625.35804933345, 
    2160.45985076257, 
    2538, 
    2993.42043707844, 
    3065, 
    2519.71484963984, 
    3053.9472021264, 
    1826.49709846625, 
    1378.49204581068, 
    2872.21052355541, 
    2262.52395275527, 
    2661, 
    1668.03383200264, 
    3084, 
    2196, 
    2002.62774404408, 
    2252.70955914101, 
    2613.36851255027, 
    2208, 
    2521, 
    1500.47930544505, 
    2424, 
    2461.12398698268, 
    2510.80506848067, 
    2954, 
    2270.14068589225, 
    2409, 
    2383.15384593079, 
    1926.91815237976, 
    2199.97695393525, 
    2089.68310942106, 
    2768, 
    3114.98168168987, 
    1112.4965591684, 
    2334, 
    2585, 
    2242.55990551453, 
    3139, 
    1880.72303455275, 
    946.842020800025, 
    1787.04288194339, 
    2880.06961066425, 
    2932, 
    2177, 
    2797, 
    1998.68778650808, 
    2821.03289642364, 
    2635.89474654742, 
    2317.14403770429, 
    2924, 
    3070.60035902151, 
    2778, 
    3014, 
    2002.75038380909, 
    2640.34680125819, 
    2722.8719548903, 
    2704, 
    2204, 
    3162, 
    2280, 
    2505.4594946559, 
    3068, 
    2048.53039940483, 
    2662.45618410226, 
    2925, 
    2827.53616125523, 
    2921, 
    2494.08485224351, 
    3038.46542137287, 
    3113, 
    917.687433621768, 
    2272.10213004935, 
    2754.10205747048, 
    1682.17776225493, 
    3014, 
    2175.31854418766, 
    2152.74736660539, 
    2951, 
    2128.99527972512, 
    2415.58087084797, 
    2471.42987092917, 
    2388, 
    2439, 
    2629.56670235254, 
    2835, 
    2598.80402366226, 
    1857.50407423076, 
    2125.34230143851, 
    2385.4506402907, 
    2417.78339607075, 
    2971.87197579982, 
    2669.97080994407, 
    2806.0501160483, 
    1632.26878025651, 
    1245.42110366654, 
    2033.00745465637, 
    2010.73028810282, 
    1964.32375228635, 
    2894, 
    1080.10750790771, 
    1364.7569137624, 
    807.070894304745, 
    3018.22095241237, 
    1376.17228592748, 
    2434.04606738417, 
    1534.11797496198, 
    2893.54599114884, 
    2388.17093650247, 
    1851.34721339222, 
    1388.21502203641, 
    3047, 
    1933, 
    1821.17287523044, 
    3228.07843824593, 
    1465.25665319977, 
    1980.01683367001, 
    2486.94932771898, 
    2613, 
    2503.71425065511, 
    1815.04097358478, 
    3079, 
    1969.48110177796, 
    1284.17663502143, 
    1904.92594063455, 
    1117.18522632049, 
    1481.84984456945, 
    2348.92693392088, 
    2814.26733192283, 
    2846.01816324337, 
    2073.95291909717, 
    2773, 
    2067.07495948191, 
    1848.64212804539, 
    2285.86503070373, 
    3115, 
    2631.24031421251, 
    2176.94879365949, 
    1522.10417398477, 
    2305.45113951426, 
    2457.05681244032, 
    2930, 
    2300.46341858479, 
    1495.85525366494, 
    804.718097058507, 
    1501.92687065495, 
    2297.86292081416, 
    2920.14938475013, 
    1370.15714132308, 
    1859.62653949662, 
    2540.79583428649, 
    2011.74261032568, 
    1857.93109127354, 
    2646.06732675923, 
    2792, 
    2642.31431081323, 
    2955, 
    2700.30226309346, 
    2552, 
    1438.45824643735, 
    1972.5281439818, 
    3018, 
    1582.71886833353, 
    2215, 
    2524.66319493237, 
    3140, 
    2032.94271060628, 
    1921.26292499368, 
    1337.83216557836, 
    1896.09010396326, 
    2584.6352170387, 
    2586, 
    3003, 
    2775, 
    1753.35590652092, 
    2529, 
    2484, 
    2797, 
    2284.2927664306, 
    2690, 
    1980.38687405418, 
    1868.49272874052, 
    1401.00818093611, 
    2061, 
    2258.11412072109, 
    2001.45470076597, 
    2186.0597336186, 
    2497.31993068393, 
    3212.92911131091, 
    1830.96870198863, 
    1790.36462311061, 
    2930.55470425278, 
    2923, 
    2618, 
    2210, 
    1876.94568028023, 
    2438.06381602626, 
    2489.94521727094, 
    2336.91067224935, 
    2276.38293538033, 
    2213.2811590476, 
    2939.73215475324, 
    1512.467068033, 
    2715, 
    2323.71688311763, 
    1982.97325094473, 
    2216.46250458526, 
    2176, 
    2836, 
    1139.01196528828, 
    2665.19155584329, 
    2535.20285019392, 
    2295, 
    1402.79799257864, 
    2575.84762366986, 
    1760.91226353329, 
    2366.54424845139, 
    1779.4440313289, 
    2568.24575142248, 
    2750, 
    2680, 
    2952.06719039184, 
    2461.49124992203, 
    2311.76872348063, 
    1570.1706164619, 
    2191.86135639589, 
    2830, 
    1991.86608249035, 
    2938.83458934059, 
    2937, 
    1208.66273770263, 
    1783.50421652516, 
    2123.640010948, 
    2049.17717358214, 
    2168.68989089139, 
    1854.86315624801, 
    2957.40727249376, 
    2360.9210780374, 
    2652, 
    2615, 
    588.219256196355, 
    2811, 
    2931.98279073575, 
    2367.09231623302, 
    1812.67047404034, 
    2592.20084591494, 
    2727.89231644785, 
    2832.00049601675, 
    1627.44185443928, 
    2274, 
    2466.21195443447, 
    1656.96558583355, 
    1383.42954633382, 
    1748.02861656777, 
    2301.64066593167, 
    2744, 
    3241, 
    2818.87351009904, 
    2153.98877328102, 
    2309, 
    3064.61439677337, 
    2116.79522340177, 
    1627, 
    3181.61928421547, 
    1658, 
    1563.51336247688, 
    2598.90205615776, 
    2670, 
    2485, 
    3079.52132739792, 
    2917.97978650397, 
    1823.19897255789, 
    3143, 
    3155, 
    2308.64538720035, 
    2592.77766744574, 
    2992, 
    2293.28066361744, 
    1377.02088581303, 
    1391.44972800904, 
    2412.47430389427, 
    2549, 
    2469.15875099936, 
    2222.03071214732, 
    2674, 
    3218.03172864753, 
    3091, 
    797.469349600442, 
    2638.67666076626, 
    2612.80409605474, 
    2880, 
    1838.02134884752, 
    2995, 
    2277.66112601257, 
    2877.10967947329, 
    1903.81008634515, 
    2098.81992783798, 
    2446.9022359541, 
    1420.26104915883, 
    2364.09741024377, 
    2510.94701832264, 
    1829.49822309454, 
    2870, 
    3183, 
    2761.22212385602, 
    2882.00834325545, 
    3032.72639679499, 
    1003.77530852664, 
    2535.31645223449, 
    1127.59587321899, 
    1372.15239477442, 
    2762.37835644673, 
    2226.9909492888, 
    2344.61090041776, 
    2092.76697636078, 
    2268.99097434785, 
    2823.30827335461, 
    1786.52227943537, 
    1726.74231073526, 
    3175, 
    2626, 
    3057.08314026789, 
    2679, 
    1662.60110014921, 
    1529.10685492726, 
    2094.16944194945, 
    1297.98432138885, 
    1546.62330931548, 
    2626.29776010873, 
    2182.28069725391, 
    1603.52749230035, 
    3146, 
    2845.84176543615, 
    2899.77275309836, 
    591.636335819485, 
    2550, 
    1871.95041612518, 
    2793.29431289756, 
    3014.19234958409, 
    3069, 
    1947.82858338442, 
    2830.07620464583, 
    2015.98473226425, 
    2510.57362663848, 
    2845, 
    2509, 
    3070.90488889947, 
    2521, 
    3056.0299950021, 
    2508.75574420008, 
    2128.69480904882, 
    2225.92619599655, 
    2879, 
    2222.13944450099, 
    2692.05524853607, 
    1894.53805337188, 
    1968.84269943717, 
    2162, 
    2221.91767712792, 
    2599, 
    2133.91134507777, 
    2554, 
    2205, 
    2457, 
    2489.66963078765, 
    2802.27446211868, 
    2361.9392415816, 
    2461.97172518644, 
    2373.2477333079, 
    1976.04562524711, 
    2262.56498665815, 
    2119.82580695233, 
    2742, 
    3224, 
    2282, 
    956.581798120973, 
    3252.83644833388, 
    1625.7426724555, 
    2789.70799896703, 
    2517, 
    2088.24986626423, 
    2882, 
    2398.48104396862, 
    2875, 
    2918.80394117152, 
    2106.66728656856, 
    2744, 
    2834.44888565006, 
    2668.23454279667, 
    2369.81772852272, 
    2414.96426013578, 
    3038, 
    2744.696403939, 
    1310.76989581187, 
    3006, 
    2021.34425220775, 
    2669.63250515323, 
    2719, 
    2716, 
    1823.62920636082, 
    3105, 
    1606.73936001095, 
    2970, 
    3106.0613447438, 
    2924.47260309425, 
    2596.03258348381, 
    3053, 
    3088, 
    2714.8861601613, 
    1144.36201374302, 
    2274.73561010414, 
    1613.52154304245, 
    3014.28627891136, 
    2186.05000083408, 
    2935, 
    2085.36156289831, 
    2413.4318877338, 
    2389.822773683, 
    2405, 
    2064.98633301885, 
    2416, 
    2822, 
    2647.38741860046, 
    1810.40560908108, 
    2357.03930340348, 
    3000, 
    1054.94168667544, 
    2672, 
    2634.47008552641, 
    1375.21963253784, 
    2070.66938741857, 
    1753.91453696536, 
    3017.8446997915, 
    816.256849375082, 
    1323.45499618479, 
    1196.91067693205, 
    2707, 
    3239.82978101457, 
    1341.96265712847, 
    2866.33451663204, 
    2070.86190885883, 
    1976, 
    3056.42197265386, 
    3070.56635718714, 
    2019.75554197626, 
    1859.2269673785, 
    1607.99630015546, 
    1536.68351501585, 
    1978.06554904616, 
    2451, 
    2556.10713780759, 
    2507, 
    3184, 
    1774.58096231019, 
    3066, 
    2056.71234923015, 
    1372.43415019134, 
    1874.11864109825, 
    1239.57530961628, 
    1727.16788031659, 
    1329.31245527601, 
    1881.5246886543, 
    1594.12960210069, 
    2792.62972278044, 
    2901, 
    2862.743690369, 
    2400, 
    2336, 
    1959, 
    2694.64230695734, 
    2257.36743639426, 
    1458.94764492666, 
    2246.99406941718, 
    2906, 
    1393.61334553503, 
    2573.59887239339, 
    1513.24051511659, 
    2820.35123801191, 
    2294.76123555673, 
    2909.53539640361, 
    2644.12987095381, 
    1404.27092538557, 
    1782.95593614287, 
    2748, 
    2630, 
    2938, 
    2701.97166526967, 
    2581, 
    1581.82654355074, 
    1903.36588756336, 
    3041, 
    1477, 
    3160.40073793457, 
    2007.85848203899, 
    1428.73230664865, 
    1955.90857409741, 
    3010.02250543471, 
    2616.19529513468, 
    2551, 
    2809, 
    2143, 
    2529, 
    1826.67370135772, 
    2059.5698796795, 
    2443.08146148668, 
    2775.6515835545, 
    2274.07536663354, 
    2735.95952166082, 
    1934.98054465941, 
    2571, 
    1266.00904830604, 
    1541.25831134749, 
    2070, 
    2460.22839611788, 
    1941.58194444746, 
    2162, 
    2855, 
    1544.37599659298, 
    2495.36342481555, 
    1627.38402708277, 
    1731.08028911247, 
    2918.16618726686, 
    2651, 
    2150.29036227408, 
    2528.47788170853, 
    2384, 
    2196.02723588387, 
    2971.6489584855, 
    2837.72645615685, 
    2658.02933213284, 
    2292.93709281282, 
    2964.43893469484, 
    2876, 
    1615.47871980453, 
    2663.95618134598, 
    2512.18938874569, 
    2328, 
    2252.74872034794, 
    2741, 
    2565, 
    2354.04410737338, 
    1631.98673940009, 
    1473.46383535169, 
    2742, 
    2972.59778896657, 
    2261.7074284745, 
    2676.14051048044, 
    2164, 
    2847.67436201035, 
    1986.72198556139, 
    3217, 
    2568.63351579278, 
    2088.86953898587, 
    2179.53608630193, 
    2540, 
    1926.02596932304, 
    2951, 
    2373, 
    2672, 
    2640.70859905865, 
    1566.6964632958, 
    2811, 
    2322.87520836979, 
    1867.42827547907, 
    2610.65582446875, 
    2666.10557246684, 
    2852, 
    1336.62571141565, 
    2374.27244014127, 
    3102, 
    1239.8532607135, 
    1609.59957087121, 
    2595.16845360501, 
    2287.00325351179, 
    2689.44331301074, 
    3242, 
    2856.34950337407, 
    2696, 
    2333, 
    1982, 
    2034, 
    1733.0457014516, 
    1778.30336655791, 
    1515.17141555504, 
    2468.95212641882, 
    3105.96833468073, 
    2915.60185551148, 
    3151.74935424679, 
    3165, 
    1134.33476369352, 
    2600, 
    2937.31543476861, 
    2969.95048251666, 
    2403.99276707745, 
    2327, 
    2507.27427902661, 
    2556.31703499434, 
    3223.40836613322, 
    3085, 
    2900, 
    2628.64537113508, 
    2574, 
    2744.24629983461, 
    2895, 
    1862.1297420836, 
    2977.3967513575, 
    2856.16738831033, 
    1855.05936179191, 
    2338.47020110703, 
    2427, 
    1552, 
    2119.94404904504, 
    2328.3560163465, 
    2910.71498149615, 
    3192, 
    2103, 
    2756.59245453784, 
    2850.4993198473, 
    2624.8813580666, 
    1240.70435137608, 
    1523.05512357279, 
    2205.82331842122, 
    2486.9743207305, 
    2361.52409486117, 
    2203.29418300581, 
    2159.0582260632, 
    3132, 
    968.836245493614, 
    1768.48034964701, 
    1764.3771129183, 
    781.498831084525, 
    3172, 
    1243.51472618712, 
    2614, 
    3041.31030929931, 
    1556.89476705256, 
    2065, 
    1372.60995002474, 
    2592.55232802128, 
    2233.62790737954, 
    1460.06991572072, 
    2832, 
    2869.1214341859, 
    3004, 
    1865.65916679916, 
    2524, 
    2797, 
    2918, 
    2002.92952956218, 
    1976.95281204119, 
    2412.30453174563, 
    2830, 
    1133.87039255308, 
    2479.83318073464, 
    3024, 
    2480.41900492921, 
    1295.46725282164, 
    1581.17808860186, 
    2889, 
    2182.97862350985, 
    2717.26207502452, 
    1942.71945661646, 
    1914.06854769199, 
    2119, 
    2280, 
    2197.15232452968, 
    2095, 
    2581, 
    2179, 
    2897, 
    2477.40309886971, 
    2477.286811612, 
    2345.77279135449, 
    2507, 
    2364.94109441321, 
    2157, 
    3024.19331220583, 
    3249, 
    2223.64085349456, 
    302.060475731854, 
    2504, 
    1934.56310961, 
    1171.14915958248, 
    3230.19121702691, 
    1736.80265650314, 
    2544.95118470458, 
    2164.9490191591, 
    2901.29459948501, 
    2357, 
    2832.95931349569, 
    2908, 
    2080.94652411827, 
    2714, 
    2371, 
    2834.15589755679, 
    2684, 
    2412.16550766717, 
    2402, 
    2990, 
    2713, 
    1432.28903156903, 
    2989, 
    2070.58301900594, 
    2715.60196216464, 
    2726.93303979032, 
    1885.55326797269, 
    2425.04387322231, 
    2997, 
    2184, 
    2655, 
    1812.09380443963, 
    2962.28140629207, 
    3090.03258156675, 
    2926, 
    3056.44497863143, 
    2837.55641221417, 
    1328.97730023884, 
    2258.44012505764, 
    3022.99408563711, 
    2221.00420094219, 
    2922, 
    2040.09319889207, 
    2439, 
    2408.79933291008, 
    2082.79088107816, 
    2379.14124022459, 
    2790, 
    2681, 
    2437.05771970067, 
    3027.45459145804, 
    1162.01411027074, 
    2674.98687385984, 
    1481.98712280161, 
    1423.65814374821, 
    2111.99620949135, 
    1810.02744937094, 
    1613.04504244543, 
    1403.98069427787, 
    2615.57205938297, 
    3238, 
    2847.99479472819, 
    1190.78006748068, 
    2037.37816471764, 
    3027.28067931872, 
    3091, 
    2092.24087941436, 
    1906.7603038311, 
    1905.34740631887, 
    1627.11036046515, 
    2010.41847515646, 
    2533, 
    2505.46940400351, 
    2517, 
    3180, 
    2131.13962074356, 
    1449, 
    1824.04725600822, 
    1785.16837683777, 
    1221.2228447809, 
    2156.54942492408, 
    2775.62705406372, 
    2182.05037728361, 
    2833, 
    2391, 
    3067.50184398971, 
    1900.0117719164, 
    2683.20624179857, 
    1358.52406268556, 
    2527, 
    2191.89822012722, 
    2880.89135580209, 
    1363.9045360417, 
    2798.59556823515, 
    2295.06319447957, 
    2709.59604373757, 
    2186.27987883038, 
    1464.70958767243, 
    1642.88543079594, 
    1664.64353318875, 
    2242.15174705837, 
    3158.32022669363, 
    2720, 
    2633.81917366082, 
    2915, 
    2744.79219727249, 
    2609, 
    1650.17289943462, 
    3064.27656719602, 
    1322.05651239564, 
    2584.58240781585, 
    3175, 
    1974.14172993281, 
    2665.14216999694, 
    2515, 
    2840.21365547284, 
    2101.9697768323, 
    2015.58004308838, 
    2795, 
    2763.98757368659, 
    1870.16885084245, 
    2613, 
    1546.2787553338, 
    2088.72291935759, 
    2504.6399792003, 
    2128.72183486287, 
    2860.04843775734, 
    1729.38441386708, 
    2385, 
    2910, 
    2682, 
    2180.07114255329, 
    1451.21086149163, 
    2560.0051566675, 
    1444.72225152134, 
    2174, 
    2040.65659079573, 
    2839, 
    2615, 
    2256.78901989155, 
    1954.97302059799, 
    2963.76401894237, 
    2909, 
    2650.8408889965, 
    2860.994173004, 
    2549.02861901681, 
    2250.02128826485, 
    1768.03926465848, 
    2728.8289216173, 
    2362.1732038092, 
    1524.54323610522, 
    2804.79990421597, 
    2986.99057885253, 
    1520.81666440905, 
    2058.75416552397, 
    3000.65233830616, 
    2867, 
    1994, 
    2862.01435812848, 
    2654.7232799129, 
    1362.52910630609, 
    2129.67866061995, 
    2196.37881630974, 
    2502, 
    2031.59608896469, 
    2938.9211805284, 
    2669.06442387661, 
    1511.32115739758, 
    2828.90321577186, 
    1667.70851976047, 
    1885, 
    2820, 
    2547.67370792761, 
    2209, 
    3084, 
    1399.5482894599, 
    1143.32917065971, 
    2624.09307141333, 
    2371.73506372833, 
    2645, 
    3226.34923270867, 
    2366.02113959687, 
    1710.15868849205, 
    1890.82664450153, 
    1947.59573512789, 
    1834, 
    1878, 
    3027, 
    2919.21815172831, 
    2144.45500579321, 
    3180, 
    1153.3006371099, 
    2961, 
    2949, 
    2843.86017238099, 
    938.842936367035, 
    2447.95315176073, 
    2567.91034725538, 
    1180.30641706691, 
    3212, 
    3224.35860377767, 
    2611.22538900308, 
    2536.42861298039, 
    2920.50527453766, 
    1883.77100135372, 
    2951.57868692235, 
    2834, 
    1816.68047893001, 
    2445.7235264299, 
    1264.09242851537, 
    2294.13846484154, 
    1547.73776030316, 
    2941.91517843176, 
    2085, 
    2746, 
    2824.44778746357, 
    1790.79413942018, 
    371.480280669141, 
    1647.5826651958, 
    2191, 
    1683.78575841916, 
    2395.00122976865, 
    2248.93419539503, 
    3113, 
    1781.70923000848, 
    2677, 
    1178.29610219977, 
    2598, 
    3229.94220496427, 
    1609.4066902874, 
    2046.60051237925, 
    1538.48811108797, 
    2554.95954995594, 
    2288.77353038013, 
    1284.04866711839, 
    3133.49708957962, 
    2814.90215591101, 
    2584.09809009499, 
    2970.94932612379, 
    1738.82012591861, 
    1216.22148894058, 
    2751.27440051577, 
    2936, 
    1920.15773097337, 
    2815, 
    2378.9045381211, 
    2447.39686285385, 
    2957, 
    3031, 
    2440.59299021032, 
    2307.95307287921, 
    1785.28972562603, 
    2946.00477114305, 
    967.613401732449, 
    1990.31391115508, 
    1848.09468605312, 
    1969.84651895182, 
    3014, 
    2169, 
    2619.32854428779, 
    2017.78874915176, 
    2148.14437394523, 
    2509, 
    2438.11840858402, 
    1346.15878795371, 
    2346.43548997511, 
    2327.82003445223, 
    2954.58158450871, 
    3266, 
    2171.32028382233, 
    2471.54850288746, 
    1896.40927787437, 
    1258.80176821875, 
    2540.31709001208, 
    3103, 
    2353.5116244959, 
    1302.6755421745, 
    2298.47471471778, 
    2073.94839185326, 
    1694.57200666645, 
    1514.92356651993, 
    2895.70403153463, 
    2052.25206035854, 
    2651.02379787737, 
    2382.77478958954, 
    2708, 
    2467.99991442636, 
    2480.84532940609, 
    2828, 
    2683, 
    1578.92709778426, 
    2989.35672749002, 
    2720, 
    2734, 
    2292.32457995472, 
    1973.15163937727, 
    1502.6088414217, 
    2169, 
    2685.97370667457, 
    2083.85182098647, 
    2914.12242644043, 
    3074, 
    2929, 
    3032, 
    2067.76356072371, 
    1394.92701695411, 
    2246, 
    2731, 
    2081.33885487636, 
    3010.29350679769, 
    2250, 
    2907, 
    2946.3298506261, 
    2448.65812315138, 
    2134.46783709907, 
    2419.79213009327, 
    2362.08122829491, 
    2764.60652963564, 
    2299, 
    2333.39108892312, 
    3055.20784849589, 
    1301.91186617553, 
    2679.73677914209, 
    2069.84092565207, 
    1784.87264985881, 
    1573.66966911775, 
    1526.16900272096, 
    1623.59490376555, 
    1868.62187008482, 
    1243.26961656077, 
    1909.012281595, 
    2180.16590666544, 
    2540.63979342976, 
    2837.66679472808, 
    2006.00332451803, 
    3020, 
    3110.40417736247, 
    2148.89097893354, 
    1947, 
    1762.933290066, 
    3225.93056675795, 
    2483, 
    2460.32892882882, 
    3175, 
    1689.8010319141, 
    2161.00680842943, 
    1561, 
    2350.20982921667, 
    2724.93340305932, 
    1855.17685651454, 
    1115.63071133864, 
    2303.7175195727, 
    2570.06219106028, 
    2424.91017829705, 
    3030.65290235233, 
    1823.88041102027, 
    1354.24909381557, 
    2558, 
    2147.12738387602, 
    1131.80267884667, 
    1232.18840955051, 
    2766.93374767098, 
    1638.40987019523, 
    2154.10396915163, 
    1487.41542828165, 
    1525.31471046625, 
    2562.23273261743, 
    2760.48519346779, 
    2001.98650994795, 
    3173.0755771154, 
    2634.20350409105, 
    2751.61273099565, 
    2638.99248685838, 
    3084, 
    1188.93551176474, 
    2325.43128621513, 
    3193, 
    1999.61494622252, 
    2854, 
    2724.03000739515, 
    2475, 
    3098.68640953552, 
    2860.22147690197, 
    2357, 
    1302.5090727689, 
    2788, 
    2510.33440088322, 
    1693.80525031131, 
    2109.89766652112, 
    2095.95699655622, 
    2875, 
    2478, 
    3233.39813849438, 
    2901, 
    2656, 
    2236.04851316612, 
    1784.71045385763, 
    2446.23985995148, 
    2598, 
    2153.54511987952, 
    2985.82894347816, 
    1633.16835501218, 
    1918.04959153929, 
    2561.8382247442, 
    2050.47858927211, 
    2464.57943455001, 
    2968, 
    1960.36983103608, 
    1401.42894739629, 
    2817, 
    2418.11319387142, 
    2709, 
    2673.73130158082, 
    1674.64790448323, 
    1501.20306273046, 
    3061.38180053394, 
    2787.57758911342, 
    2978.06393676666, 
    2835.28439778775, 
    1657.48331455002, 
    2332.02135861769, 
    2828.0429603598, 
    2863, 
    1270.12596257914, 
    2641, 
    2738.25173942838, 
    2158.23476820881, 
    2201.96939835803, 
    2473.19679654063, 
    2297, 
    2935, 
    3003.71548339352, 
    2417.75286908379, 
    2695.58250219569, 
    1430.6246794552, 
    2871.59538552455, 
    2089.61442675387, 
    2812.4711850312, 
    3068.59338364582, 
    1141.38958297141, 
    2617.25237344606, 
    1502.48568326729, 
    2293.39327342931, 
    2404.97496091553, 
    1909.88819020869, 
    1919, 
    1942.19617738001, 
    1787.12370888089, 
    2256.4537966045, 
    2759, 
    2085.62055513458, 
    1616.65883056512, 
    2944, 
    3108.18210315698, 
    1586.94608746286, 
    2640.95509930254, 
    529.588471105184, 
    2708, 
    3196, 
    2909.74320055841, 
    2135.69813822459, 
    3247, 
    2598.42100826488, 
    2506.13988011729, 
    2935.7395680525, 
    1531.02386177391, 
    2939.17044250792, 
    2371.71753765405, 
    2767, 
    1780.30398031296, 
    1497.37059668299, 
    1281.54319156615, 
    2144.62451718491, 
    2256, 
    2937, 
    2222.22366141435, 
    2751.33311418126, 
    2798.80341283451, 
    1799.53034878632, 
    1920.08344257999, 
    1688.02262110821, 
    912.053051079182, 
    2732.23248014636, 
    1615.54442220987, 
    2843.33483824381, 
    1038.34828167224, 
    3258, 
    2371.14455767024, 
    3115.83419288241, 
    3086, 
    844.172826706713, 
    1926.74249755545, 
    2709.12806690319, 
    2582.3451425001, 
    3186, 
    1655.4705732162, 
    2015.40928900571, 
    993.292703991266, 
    2518, 
    1223.13136128859, 
    1096.95255439735, 
    3138, 
    2787, 
    2581.28529622014, 
    2980, 
    2853.63443586093, 
    1914.07563797652, 
    2957, 
    2878.40579485455, 
    2292.24134672874, 
    2194.79616632239, 
    1785.47152100136, 
    2274.53148192838, 
    2414.9406295168, 
    2955, 
    3039.70721000973, 
    2411.51161407553, 
    1589.63251614951, 
    2665.52171883078, 
    1022.27351584274, 
    2019.05750268496, 
    2583.02967599031, 
    2455.75014456996, 
    2714.81587109436, 
    1936.82489336434, 
    2897.06572016693, 
    2529.73062209221, 
    2433.39214113218, 
    2420.6865305163, 
    3113, 
    2336, 
    2310.30311872561, 
    2112.9996977833, 
    2435.94844234244, 
    1694.13156067813, 
    3082, 
    2366.60715008221, 
    2560, 
    2776, 
    2023.31987029663, 
    2601.12143350597, 
    2472, 
    2432.29943083703, 
    2649, 
    1744.44983725337, 
    2998.07315175745, 
    2713, 
    2048.79839833654, 
    2708, 
    2138, 
    3057.25054614243, 
    2945.69365401042, 
    2463.21641648228, 
    3087, 
    3011.53880870348, 
    1447.99202724284, 
    2714, 
    2127.15723699879, 
    1968, 
    2284.5290271802, 
    2892, 
    2470, 
    2414.65909121397, 
    2018, 
    2340.01352348157, 
    2730, 
    2359.02289984098, 
    3082, 
    1062.67043629889, 
    1609.35775525588, 
    1929.54417338933, 
    3040.62668784262, 
    2477.05531157569, 
    2110.85605161615, 
    2841, 
    1994.07433179653, 
    3130, 
    2203.30322985344, 
    1696, 
    2435.61588527085, 
    2952.56409990843, 
    3163, 
    2219.00326527672, 
    2366.26412116344, 
    877.946936717325, 
    1758.00768355414, 
    1205.82531508918, 
    2414.89558746497, 
    1458.43355527156, 
    1514.88649985444, 
    2592, 
    2834, 
    1064.59731308374, 
    1880.64396769323, 
    2550.78316431044, 
    2195.00876569788, 
    1494.33515999932, 
    1381.98590239039, 
    2433.42650336651, 
    2743, 
    3193.80183129883, 
    2638, 
    2871, 
    2669, 
    1040.30925606562, 
    3211, 
    2012, 
    2781, 
    2436.79456758534, 
    2729.38081796909, 
    1801.99678367276, 
    2927, 
    2308.38173694, 
    2433.11812183091, 
    2118, 
    2749.65411218714, 
    2054.91594709858, 
    2872.00978727362, 
    3242, 
    1033.64915904229, 
    1213.12199367286, 
    2313.38162944663, 
    2882.99384847831, 
    2289, 
    1807.18830765211, 
    3165, 
    3054, 
    1686.79046229421, 
    1982.99552433758, 
    2501, 
    2465, 
    2963, 
    2038.16182157218, 
    1937.85063608024, 
    1198.97349221791, 
    2075, 
    1064.52917667457, 
    2820.00179366456, 
    2595.74333070783, 
    1936, 
    2689, 
    2696, 
    1564.39441894011, 
    1414.45740962101, 
    3187, 
    3106.05592529668, 
    2778, 
    1879.16733139023, 
    2724.93153455129, 
    2512.96380392419, 
    2406.16140950351, 
    2529, 
    2156.97753011798, 
    2225, 
    2417, 
    2322.34904664311, 
    2951, 
    2516, 
    1341.1135331651, 
    2846.46332108342, 
    2147, 
    2459.31810484813, 
    2736.1995009545, 
    2317.66849564203, 
    3058, 
    2064.34856325978, 
    1780.22175219557, 
    1728.00788771794, 
    1329.18802605633, 
    2449.45537298208, 
    1903, 
    1232.95983576445, 
    2266, 
    2790.66277906079, 
    2953.5321371079, 
    2037.59645522447, 
    3147, 
    2376.579119566, 
    2922, 
    2699, 
    3179, 
    1771.96175588149, 
    3259, 
    2932.45652257011, 
    2955.58213270227, 
    2917, 
    2428, 
    2751.86439100527, 
    1726.83386387057, 
    1644.95755172423, 
    1689.83851686548, 
    2172, 
    2216.46312540088, 
    2760.16402792034, 
    1912.47029230218, 
    2073.89492239971, 
    2720.19988620535, 
    2877.56957247705, 
    1731.43702088458, 
    2420.57188557218, 
    2273.32435406629, 
    1712.92115703627, 
    2303.63803064215, 
    3119, 
    3063, 
    971.213243521604, 
    2721.844774704, 
    1525.29916255205, 
    1978.47623895465, 
    2572.0721244329, 
    1667.49101463286, 
    3181, 
    1631.52299008518, 
    1717.25195995268, 
    1173.49979117918, 
    1319.19539798785, 
    2053.05953319738, 
    3134.962039983, 
    1663.54465041536, 
    2585, 
    2258.54279127502, 
    1666.61569773698, 
    2902.93693192648, 
    1200.74213394923, 
    2167.75525696419, 
    1910, 
    3149, 
    2382, 
    2944.51528719607, 
    2692.03509933639, 
    2056, 
    2807.67494503589, 
    952.24184672174, 
    1876.39045852284, 
    2892, 
    2560.95289715966, 
    2419, 
    2432, 
    1757.80387628395, 
    968.347317790924, 
    2341, 
    1698, 
    2336.38016233425, 
    3263, 
    2046.78214649992, 
    2622.53100781808, 
    3053.81443359669, 
    2391.21728226675, 
    2545, 
    1948.11913251924, 
    2768, 
    2590, 
    2527, 
    2793.71402669084, 
    3002, 
    1828, 
    3004.80847549335, 
    2707.88643827902, 
    2717.06484188597, 
    1882.01721940133, 
    2133.8986588957, 
    2733, 
    1810.33333057699, 
    2929.06454387783, 
    2451.96328488418, 
    2702.08027753156, 
    468.199488402273, 
    2704, 
    2157, 
    1991.54101263339, 
    1923.00231699278, 
    1712.8618857138, 
    2316, 
    2980.04899220504, 
    2906, 
    2489, 
    2390.03683637623, 
    2326.96120615584, 
    1948.45066439052, 
    2269.41591647859, 
    3096, 
    2090.30712353383, 
    2718.45009022882, 
    1912.21659461201, 
    3141.42062688581, 
    1830.24213550617, 
    2860.14128793005, 
    2677.40541434755, 
    3106, 
    2255.39438562526, 
    2814, 
    3112, 
    1744.69678487711, 
    810.307139341458, 
    2739, 
    1663.80423566541, 
    2177.83140047257, 
    2320.44054550809, 
    2869, 
    2425.94727754102, 
    2112, 
    2706, 
    2366.10874079764, 
    1627.07946530307, 
    2615, 
    2804, 
    1346.23826854217, 
    1315.69968627633, 
    858.174267516977, 
    2123.15142604332, 
    2453.64448132369, 
    1456.03592963064, 
    3205.00130420602, 
    2699, 
    1549.83149251931, 
    3199, 
    3225, 
    1614.26400050836, 
    2942, 
    2802, 
    2397, 
    3054.41331477488, 
    1357, 
    2896, 
    3084, 
    2818.79026010994, 
    930.784013764339, 
    2530.00147498925, 
    2133.80504068619, 
    1834.27590497595, 
    2023.1303164987, 
    2268.71047063964, 
    3223.86492582877, 
    841.882960625103, 
    2878, 
    2306, 
    2874.66302394403, 
    2335, 
    1662.39834743319, 
    2544.73621717711, 
    3047, 
    1821.64605590201, 
    2042.70697900113, 
    2456.84116765377, 
    2495.51306152266, 
    1990, 
    2108, 
    1395.1794044081, 
    2778.99279475299, 
    2598.82350515685, 
    1123.29459992097, 
    2663, 
    1365.36035083853, 
    3270, 
    2829.4617032455, 
    2759, 
    2685.82675905966, 
    2548.88941684103, 
    2940, 
    2841, 
    111.499457511029, 
    2533.84821379599, 
    1110.05651520898, 
    1141.73484861661, 
    2370.06850038197, 
    2350, 
    2120.49993534305, 
    2832.628300984, 
    2197.40867042799, 
    2398, 
    2559.88458561998, 
    3039.26485617013, 
    2078.7814323405, 
    1753.11694251155, 
    2630.34710986195, 
    2850, 
    2398, 
    2705.00991598479, 
    2475.87614410054, 
    1956, 
    2279.73706693948, 
    2321, 
    2970, 
    2060.28366562306, 
    2213, 
    1632.15922177042, 
    2370.00084240509, 
    3002.73286349181, 
    2655.48286646117, 
    2671, 
    3253, 
    2942.08930644374, 
    2976, 
    2902.55187893223, 
    2370.01576502885, 
    816.313236442456, 
    1683.49588223465, 
    1624.75211570574, 
    2185, 
    2181, 
    1472.38554565901, 
    2192, 
    1163.14290030642, 
    2899.62445912273, 
    2447.90352502985, 
    2348, 
    2355, 
    3100.08338951131, 
    3044, 
    2745, 
    2018.8855102579, 
    2570.79912101233, 
    3150.38236955093, 
    2556.12333325555, 
    1326.13057322996, 
    1938.65511725354, 
    2605, 
    2986.22226192512, 
    2902.73792267361, 
    2892.91621213163, 
    1620.98297804713, 
    2129.26647299468, 
    1985.79452342362, 
    2354, 
    2864.45616856814, 
    1997.73266064211, 
    2725.29426636613, 
    1422.90723645991, 
    2323.86953164947, 
    1733.14497282453, 
    2751.82351924135, 
    2799.37993931678, 
    1534.82899969342, 
    1791.19921906426, 
    981.140969448956, 
    2417.97070589685, 
    2433.01702554389, 
    1728.8173435062, 
    2090.11536820818, 
    2346.2332766028, 
    2592, 
    1954.26167234888, 
    2162.62124850768, 
    2021.82669343399, 
    2550.19929724443, 
    1765, 
    2784, 
    2188.11321626939, 
    2010.72026730362, 
    2888.19846045108, 
    2743, 
    3113, 
    3014, 
    2703.42594986073, 
    2701.69705331019, 
    1678.56920123937, 
    2932.71853371576, 
    2495, 
    2753, 
    2977.08280565, 
    3005.64432582148, 
    2447.71013863952, 
    2715.00277213774, 
    1969.27554558483, 
    2694.65530340151, 
    2204.98946760635, 
    1814.04061869887, 
    2525.12770400052, 
    2351.3175704649, 
    2204.86859003471, 
    2801.78187636283, 
    1054.72991471942, 
    2222.86918939436, 
    3119.23593540254, 
    1349.02581611615, 
    2811.41662074836, 
    2227.46305183304, 
    1868.64496455352, 
    771.016492563323, 
    2149, 
    2613.93463605455, 
    904.374101673218, 
    1607.18368801762, 
    2841.50135284661, 
    2915, 
    2714.04873530726, 
    1891, 
    3127, 
    2224.57784001992, 
    3213, 
    2778, 
    1164.79599175939, 
    3133, 
    1607.43515787373, 
    919.484617278758, 
    1551.75940465109, 
    2088.1260611403, 
    2483.21301285513, 
    2896, 
    966.298251140841, 
    2671.83889373433, 
    1976, 
    2389.05418450133, 
    3146, 
    2181.95525770646, 
    2319.35516310679, 
    1697.30608967988, 
    2773.50576228987, 
    2493.22033939456, 
    2181.99201645059, 
    3212, 
    2726, 
    2775, 
    2882, 
    3202, 
    3205.90845056168, 
    2063.63250967818, 
    1588.0569598751, 
    2850, 
    2358.69204138863, 
    3027, 
    2854.18584847352, 
    2869, 
    2002.05780770332, 
    835.16234005246, 
    2893, 
    2313.95292969571, 
    2382, 
    3134, 
    3039, 
    2381.80802846253, 
    2453.37905167327, 
    1342.86116753274, 
    2056.67263939378, 
    1490.39466636785, 
    2741.98690017417, 
    2911.73204629795, 
    2635.8466320524, 
    3264, 
    3078.96893099121, 
    2819.92745293432, 
    2650.58144872939, 
    2820, 
    2064.13401723577, 
    2156.44284958393, 
    2325.53572568115, 
    2380, 
    2104.03122993048, 
    2242.84821254326, 
    2802, 
    2604.1920282043, 
    2678, 
    2329.90121754368, 
    1806.02146549836, 
    3034.67323328997, 
    2576, 
    2115.49762444499, 
    2426.75048927031, 
    2505.74704488565, 
    2968, 
    1810.00344835541, 
    1844.72878480431, 
    2506.06339834843, 
    2997, 
    2625, 
    1540.10812641952, 
    2652, 
    1173.99326615756, 
    2953, 
    3240, 
    1473.53290808416, 
    594.673487937549, 
    2885, 
    1655.68519573194, 
    1486.75759354692, 
    2150, 
    2149.1978398942, 
    3004, 
    3237.09370668034, 
    640.76232738203, 
    1873.12034475957, 
    1234.91826470929, 
    2929.35439873438, 
    1865.81638745109, 
    2428.65818576946, 
    1389.91308695198, 
    2310.3218942129, 
    2397.58233221695, 
    3018.83827095585, 
    1695.95456064892, 
    2761.02593425109, 
    2070.14582300356, 
    3123.21135405228, 
    2691.27574170946, 
    2863.99044427253, 
    2942.99933137996, 
    1463.93209739463, 
    2106.83749691973, 
    1828.4319675501, 
    2420, 
    2359.90368390231, 
    1726.05856501563, 
    2732.89673099247, 
    624.388474412737, 
    2190, 
    1496.39370287981, 
    1575.60142265955, 
    2402.37977117538, 
    2335.83337135456, 
    2564.32799396499, 
    2192.65624546347, 
    2067.6972867118, 
    1837.51376347785, 
    2784.69475703706, 
    3212, 
    2986, 
    2169.57284296571, 
    2448.09098375717, 
    2071.07229479398, 
    2721, 
    2772, 
    1539.31091138228, 
    2254.12051886171, 
    2870.64655146708, 
    2596.11983742282, 
    2873.97141994077, 
    3008, 
    3015, 
    3020.13864040638, 
    2251, 
    2696.95802318288, 
    2693, 
    2249, 
    2366.45791616937, 
    2207, 
    2768, 
    1831.61507310517, 
    3026.04620446684, 
    1874.79947067302, 
    2687.85742179755, 
    2953.61859439066, 
    2306.32704578997, 
    2817.14026126092, 
    2304.84118229665, 
    2215.48253727157, 
    2832, 
    924.859685211926, 
    2531.30285555288, 
    2614.74462510643, 
    1675.32169925724, 
    2964, 
    2194, 
    1828.26636477864, 
    1633.00477597151, 
    1687.88073566507, 
    2476, 
    2618.65889636173, 
    2991.65308316845, 
    1893.08166812025, 
    3138, 
    2193.09696537775, 
    3200, 
    2760.98977403439, 
    921.812133072865, 
    2809, 
    673.549732336185, 
    2627, 
    1465.45854999921, 
    1943.32915508786, 
    2642, 
    1636.34110934724, 
    2439.17659346353, 
    2215.00789143551, 
    2590.17889490632, 
    2801.78925612132, 
    1697.42490922199, 
    1475.76871555717, 
    2232.94925884672, 
    1440.47057139176, 
    2632.56476026015, 
    550.818324013519, 
    2149.60736683719, 
    2752, 
    2754.36477715837, 
    3201, 
    3192, 
    2945, 
    1523.16676162855, 
    2324.80155802343, 
    3104, 
    1710.89849124796, 
    2547.03318331633, 
    2806, 
    2281.03971142204, 
    1188.00922470115, 
    2741.03346986742, 
    2173.64316382293, 
    2409.57155613916, 
    1441.67809879431, 
    2889.36653142918, 
    2426, 
    1845.1877996886, 
    2495.64375345632, 
    2415.94013366073, 
    2290.32276038127, 
    2118.40232276966, 
    2589.1503998124, 
    2324.6613536509, 
    3000, 
    1816.0624055929, 
    2099.78733867786, 
    1526.82925828307, 
    1984.94387364825, 
    2806.49370053059, 
    2628.25827876042, 
    1611.36016162505, 
    3040, 
    2632.85870830077, 
    2548, 
    2185.4166000067, 
    1506.09446343224, 
    2280.35017338447, 
    2408.88089512561, 
    1778.3912135377, 
    2431.77579682744, 
    2135.8998275998, 
    1561.10996405076, 
    2233.99433448707, 
    2567.62140016993, 
    1248.69821520746, 
    1948.84477097258, 
    2220.36723024661, 
    2246.54202489548, 
    2469.67610012938, 
    2540.12012415423, 
    2960.4202718588, 
    1705.87987341421, 
    2041.46252972287, 
    2229.12289623022, 
    1444.57745756269, 
    1223.58018624965, 
    2596.53934082809, 
    2136.51091890518, 
    2843.83206045284, 
    2389.00002755803, 
    1324.38819279005, 
    2035.73663755955, 
    1581.95218047058, 
    2117.53118060311, 
    2378.09583693924, 
    2025, 
    1643.87227683834, 
    1570.59985330496, 
    2953.73423241444, 
    2257.55084876358, 
    1894.32889551287, 
    2667, 
    1748.02717254549, 
    2794, 
    2593.74762983242, 
    1808.04395108354, 
    2122.60566727506, 
    1521.64071172758, 
    3153, 
    2645.70729622974, 
    1405.20588557129, 
    2837.06467641353, 
    1707.67001936022, 
    2965.01576455916, 
    1511.03016078083, 
    2743, 
    2443.98863102949, 
    2479.73543748791, 
    2704.65792954689, 
    1644.62621418699, 
    2165, 
    1253.06745712933, 
    1649.3724824992, 
    1102.49613986362, 
    2872, 
    2529, 
    1733.42611405669, 
    2321.36104129592, 
    1781.07197192258, 
    2379, 
    2235.78714425658, 
    2231, 
    2063.01223644738, 
    1219.55423773176, 
    1840.0348246324, 
    2787.2414784881, 
    2264, 
    3205, 
    2324.93531052497, 
    2140.39097972005, 
    2693, 
    1424.99611985114, 
    2732.13479866488, 
    2841.03680662112, 
    2722, 
    3038.65273291347, 
    3028.67437498031, 
    2291.9417958869, 
    2700.49011459209, 
    2443, 
    884.628618546036, 
    1945.10795469032, 
    1565.94019742678, 
    3056.61647434242, 
    2754.96632763655, 
    2135.06364575596, 
    2670, 
    1882.56500228625, 
    2945, 
    2602.25614473775, 
    2073.80268363637, 
    2239.29286883658, 
    2864, 
    2447.94704086555, 
    2558.22823467023, 
    3140.77603564852, 
    2877.57775872114, 
    1431.26236467499, 
    2780, 
    1986.2679483206, 
    2162, 
    3143.57230451614, 
    842.313874744345, 
    1555.50600867834, 
    1455.66392739845, 
    3048.92840937409, 
    1771.42320199522, 
    1728.43862494252, 
    2256, 
    2755, 
    2778, 
    1853.01621708903, 
    2515.72584317334, 
    2607, 
    1515.31382323688, 
    2525.59800485234, 
    1612.01956411488, 
    2558.27394819407, 
    1983.46119223522, 
    2994.96001293031, 
    2211.66036708896, 
    3174, 
    2556.76472963905, 
    2338, 
    2186.52043076469, 
    2711, 
    2828.25518847564, 
    2532.98932783862, 
    1938.42475317006, 
    2467.29673293178, 
    1917.05482324921, 
    2641, 
    2416.18415776739, 
    2331.00728523881, 
    2134.05760291412, 
    2312.41881864981, 
    2540.85570309084, 
    1135.11072199194, 
    1948.97170431881, 
    2076.97861374127, 
    2570.15817783099, 
    2850.50511881766, 
    2267.77102144835, 
    1819.70427566141, 
    3115.46023808618, 
    2813, 
    2238, 
    2595.33345235518, 
    1278.96401536803, 
    2244, 
    2440, 
    1830.12701918983, 
    2442, 
    1585.8467649418, 
    1625.10661964406, 
    1908.08022931158, 
    2530.85277570259, 
    1794.14043383559, 
    2570, 
    2387.2077551766, 
    1572.80838248019, 
    2462, 
    999.836918274885, 
    2398.21623822877, 
    3022.28364627692, 
    1423.94676075536, 
    2696, 
    2483.17575339475, 
    1316.55850599881, 
    2549, 
    2125.49052839496, 
    2608.7194544357, 
    2784.02227931765, 
    2142.4134270121, 
    2832.60970480033, 
    3213, 
    3189, 
    1187.46643621788, 
    455.066247503503, 
    1876.86368339372, 
    1995.83144900921, 
    1344.06800302392, 
    1221.32266459876, 
    2198.04937207688, 
    1932.10457822413, 
    3057, 
    1702.12078314503, 
    2817.9716200407, 
    2561.19386759886, 
    1975.78128356852, 
    2078, 
    2147.61073644831, 
    2603.08275874285, 
    2970, 
    2279.7149873278, 
    2725.8799946057, 
    2790.8647499296, 
    2589.17330003935, 
    2675.08737080949, 
    2548.85389907173, 
    2188.97279090367, 
    1607.6722376227, 
    2142.58136358864, 
    1356.25260348234, 
    1966.33236433775, 
    2538.22661041182, 
    1349.38300495027, 
    2239.77346292635, 
    1828.24583004822, 
    2319.85418364843, 
    1711.24152749021, 
    2412.11472409089, 
    2186.97602577078, 
    2124.83763611516, 
    2310.54449510966, 
    2345.01193106609, 
    2495.05505420114, 
    2791, 
    1312.73579927711, 
    2766, 
    3071.34148425418, 
    3025, 
    2333, 
    2775, 
    1903.34604965785, 
    1776.10833124868, 
    3068.20418324545, 
    2506, 
    2093.77559190628, 
    1589.38115856762, 
    2147.29014869996, 
    2959, 
    2035.5912768528, 
    2319, 
    1900, 
    3134.97812147465, 
    3222.85891166588, 
    2129.1308711681, 
    3162, 
    1068.67442268999, 
    1471.36521594541, 
    1540.56014622867, 
    1900.0820402007, 
    2012.0641087364, 
    2531.18665165264, 
    1613.8857137579, 
    1971.99590387133, 
    2727, 
    1325.06402452093, 
    2741, 
    1178.45406740723, 
    2600.15289814272, 
    2106.35051205462, 
    827.310760595421, 
    2574, 
    2477.92130446974, 
    1134.11349362734, 
    2407.0016284882, 
    2913, 
    2976.82782889455, 
    2262.53425831802, 
    3038.27150861247, 
    353.552220803498, 
    1380.27935109445, 
    2581, 
    2278.82301278542, 
    2687, 
    1755.55670810161, 
    2521.45706721685, 
    2840.92233987624, 
    1978.97505818288, 
    1388.43823933917, 
    2397.29741005777, 
    2368, 
    2148.15129623076, 
    2314.43270906086, 
    1986.05607315649, 
    1925.59164244474, 
    1896.41655556284, 
    1541.00437994655, 
    1405.1486273151, 
    1384.71314600506, 
    2869.44929780386, 
    2171.65876454244, 
    3144, 
    2812, 
    2290.33676628114, 
    2483.02142153373, 
    2859.82371357212, 
    2831, 
    2599.19580389381, 
    2475, 
    1871.82855009749, 
    2816, 
    2539.52320326631, 
    1511.74239899892, 
    2341.96052784731, 
    1604.29198796684, 
    1748.84780772137, 
    2382, 
    2018.48049629494, 
    2415, 
    2000.47068903088, 
    2888.54348227213, 
    2775.10054313294, 
    2779.69301206324, 
    774.075416570888, 
    2832, 
    2761, 
    2554.13047269816, 
    1511.60218189144, 
    2945, 
    2560, 
    1985.93555941731, 
    2678.21248181573, 
    3196, 
    2239.63655917953, 
    908.148063033817, 
    2802.80419382717, 
    3252, 
    3172, 
    1914, 
    1785.30798900418, 
    1962.1311584616, 
    2151, 
    2528.85805267085, 
    1684.51290217293, 
    2965, 
    1558.79171448884, 
    2280, 
    2990.96944793165, 
    1279.17396029825, 
    2340, 
    1788.44200972058, 
    3251, 
    2041.14896686843, 
    3033, 
    2712, 
    1550.71157320816, 
    889.200282885525, 
    1812.5296843015, 
    1907.28936940341, 
    2549, 
    2176, 
    2320.76251280268, 
    1973.02569603286, 
    2249.62954671941, 
    2296, 
    2117.77903651342, 
    1692.02133543872, 
    2353, 
    2802.9779885429, 
    2219.49932961243, 
    2090.13424658807, 
    2648.57127065181, 
    2619.00201115008, 
    1992.00291364685, 
    1694.28343889366, 
    2264, 
    1575.84620068006, 
    942.651260599934, 
    3024.91495024378, 
    2155.64908884053, 
    2974, 
    2688.37736481478, 
    2897, 
    2953.38460399198, 
    2299.97365832918, 
    3123, 
    2824.06470405824, 
    2876.12338511512, 
    3221, 
    1022.99696765762, 
    2512, 
    1999.42978119907, 
    2814.01956955245, 
    2745.98254181499, 
    3207.9848395025, 
    866.015421358435, 
    2607, 
    2758.86787735483, 
    2053.25296102825, 
    1014.99978265669, 
    926.991599474856, 
    2890, 
    2441.39811750732, 
    2312, 
    1884.7006167729, 
    2026.99491401288, 
    2417, 
    1584.65957274206, 
    1624.31725752732, 
    2227.26057613505, 
    2039.39921463621, 
    1628.15488522748, 
    2660, 
    2917.5536007659, 
    3053, 
    2016.05375913059, 
    1154.22519293724, 
    2858.88985185896, 
    2759.24660117361, 
    2403, 
    1777.30257920262, 
    3246, 
    2337.70039597084, 
    2315.03213809239, 
    2316.02264152918, 
    1648.45447790124, 
    2097.05326696654, 
    2890, 
    2847.11341766469, 
    2758.52540193429, 
    2319.04220331587, 
    2507, 
    1895.11843923761, 
    2212, 
    1974, 
    2911.00085052017, 
    2406.59777437491, 
    2515, 
    2791.09028495267, 
    2763.34819380584, 
    2551, 
    2777.11565450615, 
    2702.9309467099, 
    2929, 
    2572.43564480314, 
    2157.699444797, 
    2437.32074216711, 
    3156, 
    1725.88125106124, 
    2010.74035646914, 
    2091.75627677935, 
    2657.77563211581, 
    1678.40342983676, 
    1053.41077363396, 
    3012.10786223216, 
    2451.57929504011, 
    2682.59979722729, 
    2614, 
    2495, 
    2559, 
    2585, 
    2895.89539090603, 
    2333.94743028675, 
    2832.49782610331, 
    2390, 
    3190, 
    1919.00108392744, 
    2258.56872914714, 
    2758.05558784464, 
    2213, 
    2599.39410752153, 
    2411.88612122262, 
    2697.11254828829, 
    1739.24808332576, 
    2415.98506677215, 
    2256.20356345642, 
    1559.64164965, 
    2153.00801261427, 
    1927.86069264503, 
    2879, 
    3164, 
    2838, 
    1793.06603165655, 
    2919.23449052688, 
    2003.87214219937, 
    3107.98444464947, 
    2825.81022413485, 
    1660.13649125862, 
    2069.43365693928, 
    1335.14814501505, 
    3102.00248744883, 
    3079.19493658473, 
    2696.71891074311, 
    1923.95214094469, 
    1643.67676380193, 
    3210, 
    2518, 
    931.691769302166, 
    2508, 
    2674.66622931665, 
    2424.66028152974, 
    890.962081155248, 
    2696.06120990925, 
    2485.48466148123, 
    1518.5261543895, 
    2357, 
    3047, 
    516.09516437791, 
    2787, 
    2204, 
    1870.12295908675, 
    2627.03340455354, 
    2916.25134649425, 
    1892.96075015445, 
    2373, 
    2764.47194374015, 
    2433.74231668029, 
    1285.97307272851, 
    2650, 
    2225.58710600307, 
    2802, 
    2378.6971967214, 
    2553.42743729987, 
    2869, 
    2418.04716049024, 
    2001.17234205677, 
    2791, 
    1838.49538593801, 
    2540.85468812867, 
    2984, 
    2179.29936680716, 
    1910.29251696908, 
    2506.83555755272, 
    3075, 
    2482.21757437215, 
    1296.62114049337, 
    2329.88510431907, 
    2057, 
    2799.32059234517, 
    2027.07699656025, 
    2724.55899687512, 
    2918, 
    2975.26408534318, 
    2359.02234364854, 
    1778, 
    2018.67104265358, 
    2654.8212587431, 
    2753.51236150133, 
    1002.45041629237, 
    928.097432147805, 
    2168.7615375178, 
    2047.16470928997, 
    3036, 
    1006.72788822603, 
    3062.69345033881, 
    1421.70332745021, 
    2511.51963984362, 
    2570.45540349438, 
    2907.74301892084, 
    1932.4560300202, 
    2379.07653293865, 
    1320.71689730784, 
    2237.77980381787, 
    2947, 
    2424.36704084273, 
    3178, 
    2769.87690569853, 
    2322.62029068076, 
    2452.21476134206, 
    2366, 
    1820.70366685127, 
    1424.56929864264, 
    3052, 
    2173.52082889135, 
    2167.36695275487, 
    2820, 
    1884.00646992637, 
    2880.2095629869, 
    1410.72743806156, 
    2048.9978440191, 
    3086.82320597762, 
    2152.03138141106, 
    2838, 
    1192.86683586997, 
    1575.99908605267, 
    2165.33829291256, 
    1579.74058149768, 
    3111.3725976226, 
    2862, 
    3060, 
    2296, 
    1289.94547935462, 
    2001.65479833108, 
    3203, 
    2681.08422563589, 
    2145.4521833466, 
    2361.24775637816, 
    2544, 
    2735.28101631662, 
    2372.91707826956, 
    2374.45510107816, 
    2889, 
    1225.7541693529, 
    1957.24718440942, 
    1945.13189180695, 
    1707.78824462439, 
    3010.85613017039, 
    1832, 
    2202.96323714106, 
    1932.19171779803, 
    2592.94032527008, 
    1559.47131450172, 
    2141, 
    2064, 
    3025, 
    1555.45291903529, 
    806.425047826484, 
    2461.17581725048, 
    1997.01907717032, 
    1140.21222545465, 
    889.090723798268, 
    2860, 
    1926, 
    2007.33573747377, 
    2817, 
    1598.71852584287, 
    2550, 
    505.912771811634, 
    3178, 
    3135, 
    2001.64969131683, 
    2503.27808994833, 
    2195.80183573374, 
    2673.56650181885, 
    2199.20863169924, 
    2649, 
    1462.45945600627, 
    2944.19113036908, 
    2138.90737422035, 
    1856.41895686159, 
    2882.88199982888, 
    1983.89817936184, 
    2216.39390122983, 
    2566.25592205491, 
    2492.67544520073, 
    2336.268936622, 
    2666.21737636453, 
    2073.13642117156, 
    993.119136204613, 
    3083, 
    2179.72587652865, 
    2816.29620308742, 
    2825, 
    2846, 
    1740.76421238709, 
    2220.33658699261, 
    2836.36548557277, 
    1383.45855700924, 
    1747.02592597148, 
    3126, 
    2525, 
    2876, 
    2121.63851188347, 
    2471, 
    2927.02152996788, 
    1670.98776399977, 
    1481.36230290826, 
    3040, 
    2716.86067996416, 
    2130.72428699786, 
    1628.36925554596, 
    2160.62458769307, 
    1754.32317693774, 
    2339.13112013515, 
    2272.97794839172, 
    2859.24500147797, 
    2640.82380280224, 
    2445.05314079089, 
    2598, 
    3000.79664832598, 
    2200, 
    1542.99523764441, 
    2758.07646581526, 
    3019, 
    2897.60352989847, 
    2125.67292659085, 
    2570, 
    1675.8201961606, 
    2047.27795583402, 
    3110, 
    2952, 
    2696, 
    2342, 
    2717.17698576643, 
    2702.46934821318, 
    2573.91244974791, 
    2032, 
    3221, 
    2296.25650624282, 
    2636, 
    2406.43765898952, 
    2736, 
    2450.63741797645, 
    3116.61774805759, 
    2337, 
    3064, 
    2721, 
    2913, 
    2610, 
    2713.98117797585, 
    2146, 
    2623, 
    2818.13398705543, 
    2817.69474315576, 
    2532.91159121952, 
    2391.37303077926, 
    2275.69607851736, 
    1293.97836260601, 
    2636.27535848919, 
    2065.00015037162, 
    1954.5917718982, 
    2135.78917814847, 
    2538, 
    2594, 
    1285.88366062487, 
    2387.90245783036, 
    1929.56993710888, 
    2276.20406934926, 
    2123.75035266909, 
    2668, 
    1366.65045023029, 
    2079.6469441022, 
    2723, 
    2016.16812519417, 
    2477, 
    2244.25162892117, 
    2250.04481230861, 
    2250, 
    2969, 
    2483.33684825999, 
    2287.90566999708, 
    1762.34519398789, 
    2325.95303585893, 
    580.790294155237, 
    3108.04513858898, 
    2894.99766881769, 
    2709.26822613105, 
    1613, 
    2922.4013603009, 
    1959.47537036436, 
    2898.26069324142, 
    2605, 
    2592, 
    2415.02159885787, 
    1197.70267464117, 
    2076.68374710485, 
    1524.87453930282, 
    2472.3217652914, 
    2087, 
    2468.66731639575, 
    2996.75583289418, 
    2051.74306049874, 
    2113.87017572653, 
    2077.09143827016, 
    1355.17692740841, 
    2564.17477716829, 
    2667, 
    2394.7576473821, 
    1993.0329046652, 
    2083.10652184705, 
    2405.11414078209, 
    2317.31298639204, 
    2447, 
    2398.74967846788, 
    2570, 
    1882.84185595589, 
    2406, 
    3076, 
    2173.93219709763, 
    2926.38397407493, 
    3067, 
    2440.93841970772, 
    3214, 
    2528.05937410496, 
    2366.63891414713, 
    1790.82438527874, 
    2437.56890788394, 
    2536.33104722724, 
    2040.14985292931, 
    1936.28268203393, 
    1183.20478048676, 
    680.498820189325, 
    1353.61114601302, 
    1225.48347296845, 
    2539.83255069845, 
    2508, 
    2677, 
    1581.04303493832, 
    2305.11454157772, 
    2873, 
    3096.7659592257, 
    1613.46136957177, 
    2259.55369018856, 
    2643, 
    2240.98301866971, 
    1628.18070642001, 
    2245.09890300973, 
    2565, 
    2223.32832987309, 
    2300.53031538536, 
    2522, 
    2359, 
    2123.08904475287, 
    2355.84912750131, 
    2292.94709061512, 
    1295.20017408221, 
    2744, 
    2443.61866931854, 
    2670.13546629629, 
    2515.85640930217, 
    2500.35572625846, 
    2439, 
    2487, 
    3005, 
    3084, 
    3045.16124247639, 
    3047, 
    1852.70692358893, 
    1834.58142234795, 
    3018, 
    1626.09232483846, 
    2152.4853459657, 
    2871.97747321918, 
    3062, 
    1857.49779317563, 
    2711, 
    2525, 
    2175.12746465818, 
    1549.36897052574, 
    2070.73673929655, 
    1968.21915733939, 
    2837.63407926528, 
    1893.74030085933, 
    2822, 
    2606.33646835703, 
    1148.26965302495, 
    1717.97324469312, 
    1605.01758991163, 
    2308.7341843011, 
    1532, 
    2403.50768464318, 
    2836, 
    2452, 
    3151.90769569349, 
    2683.69594137874, 
    1641.29046770077, 
    2682.93704141341, 
    3110.87383407182, 
    2509.36433850579, 
    1116.49678098639, 
    1886.21273784075, 
    2373.96521636267, 
    1655.99506975696, 
    3017, 
    1365.97812085581, 
    1753.92708155163, 
    2438.56338240947, 
    1367.88092540657, 
    2805, 
    2641, 
    2538.43929679861, 
    2593.24574175356, 
    2942.54118226307, 
    2057.09710080925, 
    3156.1640674468, 
    2155.03669370941, 
    2601.9685746347, 
    2361, 
    2128, 
    3222, 
    2552.43983633579, 
    1618.74235350925, 
    2361.78326713389, 
    2271.04916280102, 
    2743.29224481743, 
    1087.92028465407, 
    2580, 
    2611, 
    2473, 
    2323.64627982905, 
    3164.98676184223, 
    2725.0810201325, 
    1814.78114614771, 
    2989.63114104061, 
    2529, 
    2092.81371735419, 
    2129.86807582401, 
    2558.34841196418, 
    2637.89622733874, 
    2746.38300692606, 
    2497.57423863049, 
    2747, 
    2061.69087398927, 
    1946.24182484924, 
    2513, 
    2539, 
    1121.18135391052, 
    2185.54684243552, 
    2656, 
    1443.33089248961, 
    3009.5047947067, 
    2103.37895898511, 
    2758, 
    2818.14485137567, 
    2283.20436197435, 
    2254.47732314458, 
    2054.03232599728, 
    2467, 
    1783.27956696376, 
    2897, 
    3184.97922238095, 
    2861.89573284031, 
    1043.66599359752, 
    2923, 
    2837.36330269637, 
    2084.86391929018, 
    2668.82773033459, 
    2633, 
    2582, 
    2598, 
    1266.33379384517, 
    1973.58604551267, 
    1860.00373389516, 
    2635.4251005124, 
    3044.0149183213, 
    2510.14386403935, 
    2161.97710474034, 
    1114.82940433079, 
    2319.34262583047, 
    2431.52182168204, 
    2775, 
    2576.60261178064, 
    2921.02048834235, 
    2425.00427687281, 
    2260, 
    3095, 
    2475.67558898134, 
    2349.86601850856, 
    3020.57184366879, 
    1941.00555927901, 
    2714, 
    2674, 
    1917.25504432336, 
    1927.28730766736, 
    1887.81081907524, 
    1285.32869631299, 
    2365.24840647862, 
    1384.80405634058, 
    2536.26353932856, 
    1819.97174123137, 
    2147.85537327709, 
    3247.35529408051, 
    2853.80079005197, 
    2854.96917652691, 
    1792.1469100339, 
    1744, 
    2658, 
    2542, 
    1089.03268428569, 
    2369.30920948761, 
    2434.32744950684, 
    2196.22694961998, 
    2502.85243491543, 
    2334.61225951152, 
    1846.21350274201, 
    2931.59769912592, 
    3045, 
    2329.19748798315, 
    2802.92166488276, 
    2629.3208703949, 
    831.086031217545, 
    2073.27691747675, 
    2198.07952553998, 
    2471.3456862661, 
    3091, 
    3075, 
    3004, 
    1973.62391108487, 
    1257.01455870277, 
    2563, 
    1915.30573832815, 
    2484.70943516037, 
    1824.68768127578, 
    2197.20633626084, 
    2798, 
    1514.18826607751, 
    1203.55765190717, 
    2501.95370191379, 
    2942, 
    2696.88377812387, 
    2112.73831220081, 
    2671.68252650877, 
    1580.48615481754, 
    2381.99733536233, 
    2492.13537773296, 
    2352.564134011, 
    2671.71031521885, 
    1660.68779949322, 
    2471.48481897646, 
    1927, 
    1626.65076442794, 
    2991.71573993672, 
    1275.63220226967, 
    1980.45931809161, 
    2379.05029164023, 
    1679.64668801919, 
    1491.72939729681, 
    2215, 
    1897.24341344792, 
    2412.87192557725, 
    2758, 
    2181.79166145483, 
    2619.34554617663, 
    2356, 
    2978.21691876188, 
    2899, 
    2468.79319030784, 
    2693, 
    2368, 
    2792.29012003829, 
    1615.08498232, 
    1956.70851890173, 
    1567.97613698948, 
    2616.72729933802, 
    2488, 
    2627.34987836147, 
    3025.71684818827, 
    852.066694587159, 
    2796, 
    2750, 
    2309.82586091575, 
    2509.92488812085, 
    2973.74097967084, 
    2731.22193174325, 
    1867.38401572281, 
    2329.71571702902, 
    2754, 
    2498.70551137125, 
    1272.70911684395, 
    2466.48270660819, 
    2221.18638394028, 
    1795.71624453293, 
    2434, 
    2240.34231217957, 
    2922.04096643853, 
    2254.56804771591, 
    3018.99453636479, 
    2446, 
    937.310696558514, 
    2077.83204881229, 
    3266.86797160363, 
    2772, 
    2987.43056193133, 
    1478.38830628428, 
    1877.87614982593, 
    2229, 
    2413, 
    2463.91679308028, 
    2219.67113373322, 
    931.733780488273, 
    2077.79102251956, 
    1847.96819835209, 
    2493.93545670658, 
    1556.06277440597, 
    3073, 
    2176.89552511831, 
    1818.04019781522, 
    2638.97443706227, 
    2211.08786228309, 
    2852, 
    2536, 
    2524.83965999798, 
    2114, 
    2279.13439608623, 
    2492, 
    2986.3884970691, 
    2721.4334034796, 
    3063, 
    2820, 
    2793.76629435033, 
    2748, 
    1751.42289054009, 
    1654.18709287682, 
    2065.47331516745, 
    2855, 
    2535.98108703963, 
    1486.07813284532, 
    2561, 
    1616.3556474295, 
    2377, 
    2255.13467312904, 
    1707.99439482685, 
    1288.55973649244, 
    2937.9676546814, 
    1461.08421684834, 
    2639, 
    1971.42035467817, 
    2314.32501361736, 
    1638.19590990245, 
    1634.83621612449, 
    3016.76631270905, 
    2301.84134679651, 
    2817, 
    2584.90070170618, 
    1479.85665428378, 
    1311.79810380736, 
    1726.30332939935, 
    2644, 
    3073, 
    2149.56348134135, 
    1478.03439892695, 
    2308.6991319779, 
    2611, 
    2471.7645724092, 
    1769.51381388338, 
    3256, 
    1996.72960668982, 
    2226, 
    2980, 
    1625.45823699653, 
    2791, 
    2516, 
    1385.29729466, 
    2707.67259621577, 
    2137.43201775255, 
    2783.52589309503, 
    1309.31746586068, 
    1488.02084439911, 
    2356.4869860815, 
    2706.26654431284, 
    2566, 
    2645.88912593977, 
    1563.52779126501, 
    2608.44866637668, 
    2375.35300820151, 
    1881.74389950964, 
    2087.6807205235, 
    2956, 
    2087.03144610465, 
    2601.084131839, 
    1486.52112557598, 
    1396.66018656356, 
    2037.77814761169, 
    1952.89153495159, 
    2919.49283475093, 
    1824.75249196517, 
    2638.301650461, 
    2553, 
    2564, 
    2486.9789384119, 
    2209.50611890412, 
    2782.55306946008, 
    2569, 
    1661.7761792388, 
    2798.30843377365, 
    1863, 
    1660.65472250283, 
    1765.05976010627, 
    2674, 
    2438.46488654988, 
    1690.6952398323, 
    1884.46698731303, 
    2503.67220797438, 
    3048, 
    2508, 
    2481.6704304937, 
    2722, 
    2661, 
    3019.49046799209, 
    2220.77496195672, 
    2589, 
    2197.78516084083, 
    2412.96659297651, 
    2626, 
    2195.3275103478, 
    2821, 
    2203.01773010533, 
    1890.99917634035, 
    2094.11926187908, 
    1392.87314783483, 
    2278.13525045042, 
    2980.73880028637, 
    2165, 
    3261, 
    2319.60190637549, 
    2473.01811847087, 
    2851.8116498557, 
    2484.50167653838, 
    2768.39500563358, 
    967.835688565, 
    3011.87475485193, 
    1999.95626766033, 
    1934.90753170302, 
    1319.58470594848, 
    2115.31859203572, 
    3115.87755419654, 
    1692.70555864825, 
    2674, 
    2637.51738037582, 
    1867.05105711098, 
    1829.16057270503, 
    2949.84730062356, 
    2295, 
    1317.74810751206, 
    1913.06331200242, 
    2563.30250291218, 
    2582.59916213882, 
    2007.53155627047, 
    2714.02028960084, 
    2224.84989209874, 
    1773.45273645871, 
    2541, 
    2782, 
    3255, 
    1530.11028158099, 
    1382.99161891536, 
    1583.4084117792, 
    2341, 
    2136.14568294203, 
    3231, 
    2371.10837158938, 
    1908.8102187273, 
    2189, 
    2290.75078187783, 
    2934.14237802143, 
    2317.34274869228, 
    2974, 
    2937.17259357746, 
    2722, 
    2141.34183915867, 
    1763.01459059824, 
    2701.83178620525, 
    3057, 
    2798.04016751068, 
    2737.91693018052, 
    2021.34282596046, 
    2602.47802194966, 
    959.367114742665, 
    3087.08150199096, 
    3066, 
    3222, 
    2252.74499357287, 
    3135.61286367344, 
    2519.31440752083, 
    1802.68694232401, 
    1213.31203832214, 
    2754, 
    2528, 
    2391.04776874744, 
    2873.32537831342, 
    2940, 
    1373.49745745253, 
    2611, 
    2090.73392545365, 
    3057.51376313931, 
    1466.79030250268, 
    2707.28757508697, 
    1784.9994451481, 
    1979.71431793977, 
    3088.0290044613, 
    2192.12353383561, 
    2604.38548591655, 
    2329.52812010636, 
    2318, 
    2576.33824371328, 
    2641.59480276662, 
    2284.07483945424, 
    1714.63846435639, 
    1823.61500032776, 
    2363.19755707668, 
    1957.48849185065, 
    2590, 
    2508.220176519, 
    2103.51377557048, 
    2368, 
    1403.37194525314, 
    1400.0186631226, 
    2151, 
    2416.91859429348, 
    2594, 
    2669, 
    3041, 
    2592.06878772326, 
    2358.72510513876, 
    3167, 
    2276.47012351417, 
    2570.07406784909, 
    2126, 
    2620.78458366509, 
    1344.35633917729, 
    1824.68409899878, 
    2245, 
    2358, 
    1917.73207847783, 
    2716.77948887344, 
    2381, 
    2131.65363548297, 
    2316.03781986389, 
    2316, 
    1928, 
    2446.99857655993, 
    2387.02726982906, 
    2257.7043850332, 
    865.873871749164, 
    2555.11918641279, 
    2639.44046710462, 
    2553.75785868888, 
    2363.02320603828, 
    1890.79624286722, 
    1528.29448371207, 
    1727.86606238408, 
    3099, 
    1799.91453582546, 
    2221.40527348998, 
    2670.05634502275, 
    3165, 
    1043.9772251485, 
    2186.96569181029, 
    2414.47607912404, 
    2912.68951077797, 
    2297, 
    3059.99904740864, 
    1658.20973294376, 
    2938.74774829942, 
    1688.63994265372, 
    2702.30712564369, 
    2731.83333836861, 
    1688.05209604722, 
    2049.48048396307, 
    971.028029770159, 
    3024.2110783875, 
    1395, 
    2198.92896010183, 
    2815.32923094178, 
    1596.99559227022, 
    2527.72545820639, 
    1594.73327924784, 
    2270.76454438156, 
    2047, 
    1710.89604402152, 
    2073.57751635, 
    2269.00296511981, 
    3235, 
    2288, 
    2035.33239123419, 
    2648, 
    2677.73624798729, 
    863.083836393754, 
    3138.42904367126, 
    1868.28442357931, 
    1932.34039760542, 
    3109.94015962109, 
    2061.30760140248, 
    1211.46569879168, 
    2182.70559833406, 
    1240.48956236111, 
    3156.80588745345, 
    2416.93736177401, 
    1630.70876790144, 
    1526.19101535778, 
    3142, 
    2534, 
    2103.50764434677, 
    1446.07210919674, 
    3033.94486663137, 
    3093, 
    2437.93231198468, 
    2386.81270154418, 
    2668, 
    1568.68311432381, 
    1569.7501114766, 
    2901.25331064507, 
    2647.84286995704, 
    1305.55135003024, 
    2369, 
    2912.58349892295, 
    1864.24300034107, 
    1386.48521761957, 
    2420.13873294434, 
    1868.50168970331, 
    2806.25893113491, 
    1912.77130790338, 
    1576.46993398173, 
    2251.993107787, 
    1970.3785673167, 
    2038.96017927248, 
    2414, 
    2313.77381647841, 
    2094.36875875493, 
    2097.12431188853, 
    2088.98888595386, 
    2503, 
    2210.55606109953, 
    2446.72831175494, 
    1280.1043440952, 
    2410.08050735955, 
    2731.01596809484, 
    1746.33752750402, 
    1756.38405874725, 
    2737.74330639009, 
    2231.94892538389, 
    1808.68666898149, 
    2635.04795171957, 
    2654.03215216401, 
    2071.6282505119, 
    1935.17150927723, 
    1630.91813747451, 
    2513.42676520938, 
    2694, 
    2705.968797586, 
    2121.87157238008, 
    2267.82484363352, 
    1679.39693420267, 
    1510.34528919517, 
    1660, 
    2690, 
    2684.91457190807, 
    2234.48853559849, 
    1925.23634740663, 
    2598.99778619716, 
    2202.99061603364, 
    2249, 
    2438, 
    2720.59008333471, 
    2212.58561647901, 
    1909.43978650821, 
    2575.32316035575, 
    2783.55073802819, 
    2628.11796672593, 
    2836, 
    2898.5264035556, 
    2477.11656779456, 
    2586, 
    2729.93899785768, 
    2471.82865172649, 
    1603.27442610963, 
    1412.65006458042, 
    3215, 
    2604.05568468572, 
    2129.52496422732, 
    2169.4893933099, 
    2247, 
    3248.05674081814, 
    2253, 
    2813.53081441766, 
    2390.19996546038, 
    2549.62655868116, 
    2818.83849222033, 
    1732.71293067144, 
    2096.4629448063, 
    1429.93029600334, 
    2970, 
    3157.39854190463, 
    1775.04262522471, 
    3067.75753894145, 
    2307, 
    1357.9098828139, 
    3084.67975943952, 
    2539, 
    2225.83854765418, 
    3064, 
    2833.58996262273, 
    1892, 
    2663.63436837934, 
    1342.59987378519, 
    1578.76820072461, 
    2061.97465831618, 
    2502.19165665115, 
    2623.54316219057, 
    1906.03924602758, 
    3027, 
    1849, 
    2501.2793781351, 
    1896.21225984183, 
    1324.74002785094, 
    1811.08143263384, 
    2415, 
    2780.5408094394, 
    2691.22008537101, 
    2124.88061972562, 
    1529.13599479478, 
    2299, 
    2367.46793713526, 
    1389.50159523171, 
    1606.5958150023, 
    738.908725181677, 
    2101, 
    2765, 
    1186.79384319162, 
    2288, 
    3088, 
    2784.60206766496, 
    1094.95234816737, 
    2693.92290731259, 
    2491.88540376983, 
    1813.95834861187, 
    2542.09104422434, 
    2178.4830781903, 
    2726.61640994911, 
    1455.68594946366, 
    1511.95375108535, 
    2848.04820898486, 
    1387.50144858596, 
    2539.58381075507, 
    2400, 
    2493.55380646603, 
    2335, 
    2068.61801755417, 
    1666.03255242355, 
    2417, 
    2620.6148492403, 
    2229.96605104322, 
    2386, 
    2338.72839882511, 
    2913.06375038151, 
    2674, 
    3128, 
    2750.31384475048, 
    1431.20449817977, 
    2244.42428647647, 
    2979.91871305416, 
    2534.8743282111, 
    2212.22543099147, 
    2701, 
    2718.22081247808, 
    2269.91168321834, 
    1718.44231526513, 
    2480, 
    2427.85656104378, 
    2053, 
    1209.46545192822, 
    1870.81275647974, 
    2412.16174272359, 
    2871, 
    3102.74354823603, 
    2575.22858115999, 
    2434.06730576751, 
    2477, 
    2467.92670925972, 
    2636, 
    2509.15349536656, 
    2571.90516505677, 
    2348.81732432417, 
    2712, 
    2683, 
    1386.17106027396, 
    2648, 
    2411, 
    2416, 
    2340, 
    2635, 
    2558.93473924595, 
    1580.72939100971, 
    2256.70107289517, 
    1736.91447345557, 
    1798.33168691157, 
    2735, 
    2200.11386854269, 
    2353, 
    2329, 
    2286.23542074086, 
    2322.08726489043, 
    2752.01701542002, 
    2612.43041213862, 
    2627, 
    1648.16686190481, 
    2940.42648320231, 
    2263.03696457965, 
    1495.87304335053, 
    2658, 
    2197, 
    3045.73017035342, 
    1571.36187146588, 
    2393.71184741646, 
    2609, 
    2321.14550602707, 
    2249, 
    1816.82199104149, 
    1517.49091722929, 
    2742.97951047741, 
    3144, 
    2319.68467212895, 
    2428.25590014471, 
    2156.20088012021, 
    1359.48929620908, 
    1860.94478192677, 
    2842.82818923714, 
    2848.69410560891, 
    2810.99885916007, 
    2825.53269385226, 
    2388.83790765712, 
    3010, 
    2938.33755892601, 
    2952.9961700067, 
    2616, 
    2867.002582268, 
    2941.70242140932, 
    2673, 
    2633, 
    2482, 
    2364.36716040424, 
    3057.67048721935, 
    2398.56868542291, 
    1852.68738917907, 
    2124, 
    1430.97260108717, 
    2382, 
    2431, 
    2561.08932131603, 
    2457.42379210159, 
    2269.00408619679, 
    2913.59921347433, 
    2947, 
    2105.9206488062, 
    2085.74049674929, 
    2606.57044858085, 
    1939.84405241895, 
    2435.2498098741, 
    3081, 
    2174, 
    2468.68524379083, 
    2557, 
    2509.8777162863, 
    2301, 
    2294.8937737261, 
    2281, 
    2715.00200560994, 
    2723.85288945451, 
    3011.78077598286, 
    2984.67318582913, 
    1868.0258377325, 
    1005.08287966774, 
    1271.48384124285, 
    1650.85883857487, 
    1476.82953532695, 
    2457.08996439581, 
    2383.96535984589, 
    2652, 
    3124, 
    1238.03533569281, 
    2611, 
    2859, 
    2579, 
    2434.37876805124, 
    2389, 
    2505, 
    1584.64545403002, 
    2440, 
    2551.80971134055, 
    1909.71783246077, 
    2553.33773386306, 
    2392.02270889449, 
    3124, 
    1950.97366753285, 
    1368.45745439146, 
    1765.31349672041, 
    1261.23635385652, 
    2540, 
    2409.53232142503, 
    2449, 
    2664.16571258574, 
    2570.25597358223, 
    2985.32373216319, 
    2389.0344116278, 
    2385, 
    2453, 
    2516.05697977829, 
    2658, 
    538.8626293984, 
    2253.33808186584, 
    1108.22951168839, 
    1648.64340804557, 
    1167.62011005956, 
    2310, 
    2550, 
    2731, 
    2400.06128899134, 
    1519.63946863431, 
    3155.61403304178, 
    2422.96994597131, 
    2350.07132256509, 
    2629.17688034266, 
    2660, 
    1605.96110811238, 
    2780.40698759795, 
    2338, 
    2500.16923642505, 
    2244.96362529446, 
    2711.53453601187, 
    2847, 
    2137.6984856596, 
    2971.22578800201, 
    2999, 
    1923.19352542631, 
    2277.5574313832, 
    2490.04644283994, 
    2635, 
    2403.32838735133, 
    2577.4132709282, 
    1951.88347628477, 
    1346.38739265217, 
    2098.59890338923, 
    2431, 
    3019.69258709038, 
    2079.90205909083, 
    2659.32856664435, 
    1684.90327391754, 
    2426.46681210786, 
    3059.79352058445, 
    3039.47394141363, 
    2942.80340330978, 
    2544.51855170939, 
    1564.63422791783, 
    1752.61545745587, 
    2797, 
    3231, 
    2732.37506878685, 
    3032, 
    1872.5690947753, 
    1851.25254447555, 
    2914.14406622821, 
    2622, 
    2415.61173490644, 
    2387, 
    1321.90844783131, 
    2886.11803298904, 
    2373.46620678639, 
    2410.91476949235, 
    2612, 
    2482.66032231861, 
    2965.17773453349, 
    2579.02290182909, 
    2452, 
    1643.0024365213, 
    2964.92338248589, 
    3105, 
    2905.21847468991, 
    1963.55631464944, 
    2499.67680259308, 
    2317, 
    1464.5180196773, 
    2487, 
    2415, 
    2358, 
    3039.83813419699, 
    2437, 
    2984, 
    2464, 
    2387.0850350591, 
    291.005977186473, 
    175.344424818922, 
    522.20509244341, 
    691.86213585919, 
    732.127554977613, 
    799.236771715167, 
    1071.7320510743, 
    634.265135803135, 
    1222.39147949384, 
    1511.0471893712, 
    791.197868962717, 
    42.4317623463531, 
    39.4090445641522, 
    53.0086245452034, 
    1218.56134978161, 
    938.145567416382, 
    993.790287799281, 
    1708.57428068677, 
    342.894735402686, 
    984.416354022211, 
    977.093261615287, 
    1446.04109660547, 
    1980.7074702297, 
    1051.65158093215, 
    115.389218367469, 
    170.976123986414, 
    928.303329237382, 
    673.748838458329, 
    1235.95498045986, 
    611.135805897386, 
    784.653859335245, 
    1683.00888999643, 
    721.258976472161, 
    903.888781425779, 
    1226.44615316995, 
    1852.07763350216, 
    961.382143265069, 
    688.746646687673, 
    1826.90981333553, 
    785.369015198342, 
    594.435583456291, 
    1989.37764801136, 
    1416.700359402, 
    871.139676581491, 
    776.288183175935, 
    749.187053250588, 
    1183.73420289345, 
    851.944092184909, 
    182.012289117099, 
    445.059456939393, 
    428.152822232131, 
    515.083269869726, 
    740.895198228842, 
    423.08282895375, 
    2027.39102193326, 
    743.250476359854, 
    824.87805064709, 
    1149.20641584006, 
    1110.18696296175, 
    753.94255757905, 
    202.851436477279, 
    392.188301045624, 
    984.753939435826, 
    587.701421300324, 
    534.578264330353, 
    2247.60375694377, 
    1130.36910850281, 
    1242.00453076995, 
    504.885755691272, 
    292.410024453932, 
    139.34008339514, 
    730.364724966286, 
    837.013187234724, 
    1369.49705046536, 
    1098.80941689203, 
    67.8635575617012, 
    892.179751006673, 
    944.358470061781, 
    934.817167930535, 
    537.309071553093, 
    605.00997084508, 
    1345.76293855094, 
    2128.27291930599, 
    1038.15719938358, 
    1079.31396484439, 
    849.028381049462, 
    386.079659908441, 
    574.427729565641, 
    307.92785041692, 
    929.311254947315, 
    1290.56108594757, 
    54.7042936172119, 
    901.026594680972, 
    1320.63298634181, 
    1791.29254055017, 
    1914.70077054864, 
    665.750197936132, 
    588.961527086485, 
    655.541858435545, 
    586.571755628414, 
    694.999002359353, 
    920.455631797343, 
    965.406995740147, 
    956.25729865355, 
    283.456528022659, 
    400.473872518334, 
    765.331263950242, 
    654.863531518282, 
    777.749208520103, 
    1789.54228163659, 
    972.966302925052, 
    894.0301922434, 
    851.653072078683, 
    226.263296708841, 
    722.064236411112, 
    636.181260792633, 
    915.314077024057, 
    400.963156998843, 
    462.264617599467, 
    603.11108182468, 
    404.124187790032, 
    1302.31349909816, 
    718.252254405791, 
    659.695325142622, 
    1075.65697121898, 
    1574.47723482265, 
    1061.93112316708, 
    559.560925636289, 
    295.535442706836, 
    783.831514841085, 
    787.171801994776, 
    1000.92212665233, 
    444.010599009296, 
    1056.81844885358, 
    929.297053817434, 
    801.583011958587, 
    48.6544679282023, 
    331.068191425198, 
    150.204841718667, 
    408.323528914525, 
    778.853392782645, 
    973.957022278616, 
    1745.23830452214 ;
}
