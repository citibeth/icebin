netcdf _elev_mask {
dimensions:
	time = 1 ;
	x = 76 ;
	y = 141 ;
variables:
	byte mask(time, x, y) ;
		string mask:units = "" ;
		string mask:coordinates = "lat lon" ;
		string mask:flag_meanings = "ice_free_bedrock grounded_ice floating_ice ice_free_ocean" ;
		string mask:grid_mapping = "mapping" ;
		string mask:long_name = "ice-type (ice-free/grounded/floating/ocean) integer mask" ;
		string mask:pism_intent = "diagnostic" ;
		mask:flag_values = 0b, 2b, 3b, 4b ;
	double thk(time, x, y) ;
		string thk:units = "m" ;
		thk:valid_min = 0. ;
		string thk:coordinates = "lat lon" ;
		string thk:grid_mapping = "mapping" ;
		string thk:long_name = "land ice thickness" ;
		string thk:pism_intent = "model_state" ;
		string thk:standard_name = "land_ice_thickness" ;
	double topg(time, x, y) ;
		string topg:units = "m" ;
		string topg:coordinates = "lat lon" ;
		string topg:grid_mapping = "mapping" ;
		string topg:long_name = "bedrock surface elevation" ;
		string topg:pism_intent = "model_state" ;
		string topg:standard_name = "bedrock_altitude" ;
data:

 mask =
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    2, 
    4, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    2, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    2, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    0, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    4, 
    0, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    4, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    4, 
    4, 
    4, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    2, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    2, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    0, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    0, 
    0, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4,
  4, 4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    0, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 
    4, 4 ;

 thk =
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    619.76062172489, 
    659.866111713342, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    825.097509870139, 
    711.409306576301, 
    1048.06924397297, 
    944.352535799662, 
    728.399537362042, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    812.916983291322, 
    984.888866911745, 
    851.833155627868, 
    1121.48016839911, 
    1073.15000592064, 
    745.70588071795, 
    0, 
    0, 
    0, 
    0, 
    1046.10557622849, 
    817.194092008417, 
    648.104453756767, 
    496.689859553048, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1109.45156511236, 
    918.143767507366, 
    1494.4905580327, 
    914.753434514587, 
    926.715713734178, 
    791.335962058119, 
    0, 
    0, 
    0, 
    0, 
    811.569742821831, 
    826.432996164173, 
    671.717222253676, 
    720.10851106215, 
    628.201057432141, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1016.5196655638, 
    832.379081158835, 
    958.099122291247, 
    1079.98262702109, 
    1031.94298579516, 
    883.29452818003, 
    922.561336652408, 
    0, 
    0, 
    776.277993069761, 
    1021.67303195921, 
    849.154909992748, 
    1141.00745897432, 
    661.93054377379, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1114.8416189916, 
    1077.53683134373, 
    951.835055787895, 
    960.696426308658, 
    1211.21113241265, 
    1187.19239224852, 
    1032.42750730019, 
    1230.25041254444, 
    0, 
    729.417817852786, 
    774.232810691747, 
    1011.50818199045, 
    921.534460059671, 
    831.969544155846, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    40.339036854319, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1149.60545169545, 
    924.27004236242, 
    988.238353064582, 
    1393.44290684693, 
    1320.9994617514, 
    1257.74855334507, 
    1148.27333029259, 
    1092.99702048945, 
    1388.0952324981, 
    987.351432535899, 
    978.139363003669, 
    1118.84485937384, 
    881.925017680448, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    25.6979138849817, 
    768.546627224854, 
    772.80342252862, 
    1057.67444446924, 
    856.562299890687, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1230.13738569694, 
    1093.50538419547, 
    852.242902068921, 
    1230.94676377054, 
    1380.35861963468, 
    1378.86959435095, 
    1428.23705152363, 
    1356.2990061184, 
    1623.46296841114, 
    1506.84844237116, 
    1185.057007167, 
    1176.05619906781, 
    1154.80658336551, 
    960.180608787342, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1.10805892750776, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    751.367335464617, 
    674.60468603184, 
    679.222814721228, 
    961.905808781495, 
    1241.54207206463, 
    858.528635459555, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1216.07215664384, 
    1193.23893020971, 
    946.736510304772, 
    1338.53694569629, 
    1478.30404887487, 
    1478.93164033879, 
    1555.49012002273, 
    1432.49426570147, 
    1501.05604956544, 
    1393.66376875366, 
    1365.44256017554, 
    1330.41148823838, 
    1267.58338947436, 
    1183.7528471513, 
    1004.74177348306, 
    903.82845233372, 
    722.762411240928, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    915.196899385979, 
    854.986867132413, 
    937.637143902022, 
    890.051861174933, 
    854.521017705946, 
    689.984390001348, 
    0, 
    0, 
    0, 
    0, 
    828.853068120213, 
    846.109368909941, 
    0, 
    840.833954521373, 
    1160.65405974657, 
    1053.25851391938, 
    1262.43826409395, 
    785.238097202789, 
    1150.46071840991, 
    1045.43739870872, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1248.13029613876, 
    869.5100506023, 
    1472.89752189176, 
    1404.91336646428, 
    1308.36554115634, 
    1577.9755725803, 
    1638.3386402098, 
    1623.86109715914, 
    1598.72796625636, 
    1561.91446118166, 
    1557.95227520525, 
    1415.81215441987, 
    1509.34830695016, 
    1371.3378789744, 
    1298.8265570871, 
    1169.67737735787, 
    1032.07581329642, 
    895.018269660462, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    744.199876321737, 
    785.184866218496, 
    935.640474697838, 
    1009.30376863974, 
    780.205396896848, 
    849.57677365962, 
    719.664569452508, 
    760.593964827876, 
    718.969621023538, 
    783.306388631144, 
    1063.72302504637, 
    1117.44901509906, 
    939.40687243765, 
    986.140981320631, 
    1384.52658885823, 
    1292.68185506124, 
    1142.38150968619, 
    1385.68290262729, 
    1211.6417079323, 
    725.470217027374, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    850.781074985942, 
    1106.02552548622, 
    1092.90671684806, 
    1115.6675437292, 
    1140.40059688912, 
    1098.78024931457, 
    1033.78235538703, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1054.26060099517, 
    0, 
    0, 
    0, 
    1236.07076688952, 
    1175.20026914567, 
    1277.1443765334, 
    1329.96019901848, 
    1471.89889850889, 
    1556.31553124628, 
    1438.80409784012, 
    1621.05852671124, 
    1734.16960276197, 
    1782.1461281017, 
    1769.8505115922, 
    1694.71626978064, 
    1647.87799680837, 
    1571.3980963892, 
    1526.57914223212, 
    1400.76512384044, 
    1293.14383911053, 
    1159.37886000557, 
    970.370462667695, 
    788.345908772184, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    821.133714628741, 
    677.820689199461, 
    1101.66803123666, 
    725.899265899717, 
    759.072160747092, 
    848.163367295273, 
    848.975063964148, 
    861.124511114681, 
    846.085955497531, 
    770.388186993001, 
    812.070454221835, 
    973.588517226259, 
    1008.07561175581, 
    1206.15089368436, 
    1249.14497044304, 
    1416.42608615576, 
    1403.84649995531, 
    1044.13317280214, 
    919.873719460169, 
    824.433897715475, 
    805.990350167109, 
    783.336072639284, 
    769.929961487314, 
    916.930209216607, 
    857.174927817443, 
    546.092398453123, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    975.677825218322, 
    1009.74511216299, 
    0, 
    1039.80460045216, 
    1369.58463598308, 
    1351.34752256242, 
    1331.50181555014, 
    1343.48694512426, 
    1269.24884633841, 
    1251.29513096951, 
    1215.33579966039, 
    1158.72249501759, 
    1116.85139617262, 
    0, 
    1123.31220194222, 
    1627.50679630071, 
    1215.35116011277, 
    1074.86704551163, 
    1227.74402986159, 
    1334.43626583889, 
    1393.3216306963, 
    1408.02880940033, 
    1372.20279357641, 
    1596.10439056619, 
    1696.79258091442, 
    1790.02541503578, 
    1747.45001213287, 
    1797.19713036456, 
    1836.47813618452, 
    1846.80985600214, 
    1803.64142016167, 
    1776.6448019445, 
    1695.11542294163, 
    1568.88674372948, 
    1481.4401105053, 
    1370.66818280037, 
    1226.62294228785, 
    1111.31632588108, 
    1017.1106254501, 
    1095.82512336609, 
    1164.39910827571, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    859.484384435952, 
    736.166102366295, 
    981.031497988958, 
    895.472898906697, 
    936.823527769207, 
    905.066919612614, 
    902.829682781642, 
    929.480402429471, 
    1101.88852917966, 
    1073.40278424195, 
    1140.0228588005, 
    1266.70301857625, 
    1496.5246820425, 
    1598.45968629854, 
    1721.66710494163, 
    1352.732777312, 
    1052.06852285635, 
    1021.73997591339, 
    1070.70914404475, 
    916.795190043235, 
    914.398811056475, 
    1044.03196977714, 
    1052.07552696313, 
    1048.57911411558, 
    1033.86020936612, 
    816.87533466129, 
    752.776334782679, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    757.626244429693, 
    966.90659935721, 
    754.443641488614, 
    876.334702307485, 
    913.664836416339, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    718.090899897281, 
    1250.49385531175, 
    1467.64792500394, 
    1116.80727454385, 
    1247.79615091684, 
    1314.57006181027, 
    1227.49215819705, 
    1320.28055657044, 
    1240.60777013512, 
    1168.45794186993, 
    1411.83940592321, 
    1312.85731899466, 
    1265.14071895248, 
    1187.21291582059, 
    1365.17233541207, 
    1471.47703263868, 
    1376.0272032483, 
    1181.03291567189, 
    1534.54410778114, 
    1395.9979864265, 
    1578.34212290171, 
    1443.72841418352, 
    1592.31399148555, 
    1685.56738422834, 
    1705.88568720742, 
    1860.20313737261, 
    1867.30640381013, 
    2011.47048554915, 
    2032.6006147975, 
    2047.47175967335, 
    2049.19715000422, 
    2038.70718201914, 
    1841.39224790296, 
    1659.88726299352, 
    1551.82927392992, 
    1462.23794205688, 
    1368.14078249014, 
    1248.18377213524, 
    1192.6358453167, 
    1283.73054426478, 
    1232.82724980005, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    699.432137037739, 
    591.269700960831, 
    802.452919971314, 
    877.085237244409, 
    1007.78661720836, 
    1162.22534538041, 
    1131.13434728833, 
    1139.68200563708, 
    989.177189474941, 
    1250.70419903456, 
    1425.68370666393, 
    1443.68606159941, 
    1675.69476606671, 
    1297.24608821846, 
    1487.07821375595, 
    1623.42721253043, 
    1458.87294344229, 
    1468.06722900131, 
    1174.24894608844, 
    1219.43202667095, 
    1346.47494533004, 
    1323.67142461483, 
    1300.07071695785, 
    1336.40478879011, 
    1291.55635916418, 
    1304.8761988231, 
    1316.65506552782, 
    1214.74245967963, 
    928.260113033049, 
    552.182106866976, 
    695.836317995385, 
    904.834766851415, 
    829.223509874214, 
    970.102765625321, 
    813.957435471379, 
    0, 
    0, 
    834.077100876961, 
    1002.50310421598, 
    1012.79045958266, 
    1041.79390239826, 
    920.834885961522, 
    920.10249130088, 
    875.980289404084, 
    840.35751014825, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    960.307696512337, 
    1499.86061984725, 
    1482.52003044028, 
    1445.49328711123, 
    1394.5099952163, 
    1474.84349848745, 
    1465.98681832413, 
    1397.98564937342, 
    1410.95871518691, 
    1592.47128259901, 
    1401.82023675545, 
    1392.64921329653, 
    1448.11657687603, 
    1427.97441717398, 
    1587.13335276044, 
    1404.18468034047, 
    1477.20046189174, 
    1356.89552954405, 
    1337.26133670914, 
    1581.08218311153, 
    1584.07992494084, 
    1643.53480134764, 
    1839.9135172624, 
    1839.01369186528, 
    1731.82649626549, 
    1892.58166096057, 
    2067.48536094475, 
    2208.49686918768, 
    2307.99379568281, 
    2289.52300996983, 
    2205.98166998878, 
    2006.85376951579, 
    1841.61163610106, 
    1731.8873438043, 
    1625.0524902678, 
    1581.79396050998, 
    1495.33725601124, 
    1406.14374697054, 
    1384.90848052318, 
    1395.73431539946, 
    1389.50809012698, 
    1312.66042973395, 
    1138.63662181227, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    647.28964499849, 
    721.190419708062, 
    908.792026840252, 
    1097.71050333435, 
    1329.96543409664, 
    1571.56425380684, 
    1504.02718840732, 
    1266.88813048795, 
    1405.60954057213, 
    1553.02584788115, 
    1802.58665573467, 
    1718.49791403217, 
    1687.77664655807, 
    1556.23028968179, 
    1621.33623874828, 
    1837.12632263595, 
    1907.66319047474, 
    1773.80354402758, 
    1519.82464057613, 
    1516.35393294492, 
    1663.28692822183, 
    1675.10327920522, 
    1591.40214754922, 
    1609.04391259742, 
    1473.48768853987, 
    1424.53087594193, 
    1345.86375686575, 
    1247.98870878533, 
    1054.42802536241, 
    955.108010744325, 
    949.324418407881, 
    987.287241513439, 
    1102.05966226112, 
    1251.89325514544, 
    1068.00555658401, 
    798.917214370981, 
    818.369969275709, 
    936.435356812067, 
    974.166915237533, 
    962.134682315935, 
    1066.35818467849, 
    1037.19361153591, 
    1054.51776079927, 
    1117.34300567623, 
    1105.43848669866, 
    0, 
    700.821568922845, 
    1012.32519725862, 
    0, 
    959.70810730934, 
    977.092060782394, 
    0, 
    0, 
    0, 
    0, 
    1005.88662976217, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    555.759090591934, 
    743.888055807307, 
    1072.66842211043, 
    1429.30738855329, 
    1382.85348135596, 
    1448.58769554641, 
    1578.98383340249, 
    1632.53772513707, 
    1804.29935432004, 
    1689.26247052283, 
    1673.19817320087, 
    1637.80677973013, 
    1413.71544054283, 
    1434.52997542808, 
    1503.78165755636, 
    1534.09181173412, 
    1528.11857615531, 
    1518.40522892954, 
    1588.84156561304, 
    1509.96872405518, 
    1480.26244356056, 
    1623.8101645493, 
    1675.21840699032, 
    1706.36607131473, 
    1754.49868827346, 
    1995.22960267547, 
    1949.08017707865, 
    2056.18276825169, 
    2197.93298216972, 
    2299.96450689612, 
    2437.49381671306, 
    2356.04428573041, 
    2031.91157624305, 
    1922.26384081089, 
    1921.70734120405, 
    1867.17557322243, 
    1782.25600489922, 
    1706.37074862821, 
    1609.08445973635, 
    1525.56541207646, 
    1534.29953071102, 
    1571.13505736105, 
    1513.5103900698, 
    1618.06952604953, 
    1175.26276287732, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    689.656661148165, 
    0, 
    0, 
    0, 
    789.530291423017, 
    965.72076274162, 
    1135.41391098644, 
    1462.07200541843, 
    1615.80291211628, 
    1723.8612643952, 
    1672.58733655465, 
    1417.13124764588, 
    1456.41154177587, 
    1774.86612621583, 
    1862.27159342229, 
    1839.58332752937, 
    1776.74762431996, 
    1796.00646462973, 
    1845.32260190769, 
    2027.07687130049, 
    2034.50154911068, 
    1833.41923157532, 
    1678.40059156818, 
    1608.22051165521, 
    1508.4371283612, 
    1604.49954405539, 
    1711.20391193285, 
    1618.56715373021, 
    1552.28720010653, 
    1582.46406750776, 
    1522.20167400104, 
    1437.15053453036, 
    1258.40633353684, 
    1084.44390382312, 
    1093.59636659233, 
    1254.5462236326, 
    1335.32229663567, 
    1426.24892998542, 
    1302.40056307256, 
    1080.72812248474, 
    1053.04002682002, 
    1052.96832548951, 
    1130.94614299971, 
    1137.64676017196, 
    1272.99676082051, 
    1506.25726865132, 
    1393.54115734846, 
    1301.09603469609, 
    1072.60191770635, 
    1632.21112458646, 
    1528.03424885193, 
    1057.84580956466, 
    1108.08032754758, 
    1256.67990412834, 
    1275.817693471, 
    837.998042854568, 
    1248.21089311493, 
    1286.20187269529, 
    0, 
    894.995592107849, 
    1167.87508275357, 
    989.489567394933, 
    1595.45388697459, 
    1076.48728412698, 
    488.02040064753, 
    844.978264823533, 
    475.277009098289, 
    1047.10126038692, 
    984.75745357399, 
    1348.36196688427, 
    1495.86284333289, 
    1616.09069281734, 
    1599.08934544199, 
    1603.30964430853, 
    1582.70511318366, 
    1682.70162880783, 
    1741.44095323814, 
    1771.34717089638, 
    1772.43738988446, 
    1725.92210442383, 
    1643.79658585467, 
    1714.07973186909, 
    1572.63675314631, 
    1501.07475078586, 
    1527.02086921968, 
    1594.23605142846, 
    1499.45921465781, 
    1444.88174730666, 
    1597.80106217578, 
    1637.1291025901, 
    1932.8890046902, 
    1926.31750406338, 
    2113.29392997716, 
    2193.689459322, 
    2311.98838023582, 
    2320.07545365322, 
    2463.76100974861, 
    2434.87822112836, 
    2221.95972719127, 
    2096.00771361791, 
    2095.93562156619, 
    2159.52957166078, 
    2041.54774668138, 
    1925.14559726757, 
    1862.9086628531, 
    1739.89928964545, 
    1673.57277819735, 
    1624.21537782728, 
    1610.32411912292, 
    1567.90723629264, 
    1511.02103626361, 
    904.346031857671, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    789.858354070739, 
    946.787174878334, 
    662.998505977, 
    560.446978400459, 
    917.117684018133, 
    1114.84735825345, 
    1414.28048212707, 
    1579.93441858417, 
    1621.00786752169, 
    1700.9060177844, 
    1730.06023253091, 
    1610.03715438601, 
    1484.89506879941, 
    1739.89500014405, 
    1981.36917035713, 
    1895.35307375409, 
    1868.13450674869, 
    1975.45353983308, 
    1964.95306752245, 
    2190.44694518682, 
    2132.78504438448, 
    1921.39102838394, 
    1854.44505697771, 
    1809.3861197238, 
    1663.51021414897, 
    1584.79091195112, 
    1713.6734815088, 
    1620.7960041647, 
    1661.12414397797, 
    1757.78747900461, 
    1686.75262726525, 
    1534.13455807889, 
    1369.48220694643, 
    1232.62382540196, 
    1276.69750071673, 
    1429.74628452219, 
    1447.05665696168, 
    1426.95957443829, 
    1454.86553334129, 
    1341.60122636642, 
    1367.61084159812, 
    1368.52352486711, 
    1346.16068615101, 
    1456.41024159405, 
    1574.68788251934, 
    1729.56219709911, 
    1511.32684362544, 
    1340.92516904907, 
    1487.38985116874, 
    1526.5562148319, 
    1344.90303033412, 
    1239.23896356904, 
    1250.14416361309, 
    1352.25739506263, 
    1334.55949510341, 
    1151.58628690492, 
    1301.93226056424, 
    1120.85757306815, 
    1164.12836160518, 
    1022.35724309709, 
    1000.94870920042, 
    1304.05918363494, 
    917.72526479195, 
    1019.34707910172, 
    1841.82309299182, 
    1083.79337316215, 
    1109.67129802193, 
    1348.17776112675, 
    1360.04023636377, 
    1443.20614510634, 
    1657.54812050667, 
    1749.94238850374, 
    1737.73632848912, 
    1692.029350006, 
    1644.83738052979, 
    1624.59835050182, 
    1702.67831292052, 
    1802.9852366731, 
    1773.97492735799, 
    1647.60004198163, 
    1653.79533870586, 
    1591.23348484796, 
    1550.56131681892, 
    1536.20576013036, 
    1604.19550174649, 
    1595.05644540977, 
    1776.43473750868, 
    1561.96892344327, 
    1605.35716437198, 
    1728.11962263038, 
    2072.28512416464, 
    2248.39130543967, 
    2196.81357847634, 
    2217.51641719219, 
    2426.78247022116, 
    2447.31283980884, 
    2471.53639428403, 
    2369.94741305126, 
    2272.69208566771, 
    2234.10720307467, 
    2227.96908537598, 
    2269.54149544049, 
    2083.5912612554, 
    1970.66850011234, 
    1986.52898791977, 
    1866.09427637214, 
    1759.79163785712, 
    1709.12943051821, 
    1650.12726137819, 
    1623.09552256218, 
    1176.94427192887, 
    902.31689030284, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    777.310668255752, 
    826.397534546392, 
    1166.61241410147, 
    975.97767389774, 
    906.941745905761, 
    775.162149290472, 
    1050.15577387961, 
    1222.25379016456, 
    1443.38605584548, 
    1422.38995169385, 
    1537.66426559915, 
    1806.49690650068, 
    1897.10738823708, 
    1709.5982002957, 
    1666.40663681552, 
    1569.68948899279, 
    1746.91981570139, 
    2019.25620086298, 
    2132.76673955925, 
    2141.77742437619, 
    2159.62205508093, 
    2239.95506163701, 
    2219.11232120041, 
    1990.46840409255, 
    2034.85904839755, 
    2003.55643463658, 
    1817.83655528453, 
    1731.47371150791, 
    1732.81462847488, 
    1663.26587429391, 
    1727.58059093793, 
    1753.94809599643, 
    1655.2271443023, 
    1566.50327455796, 
    1443.49506383011, 
    1515.04812696158, 
    1578.38521399729, 
    1633.85292086788, 
    1586.92336201532, 
    1493.76855496376, 
    1500.95007887109, 
    1592.55147936146, 
    1649.49786102945, 
    1635.66188983127, 
    1752.94209649327, 
    1630.05363359034, 
    1664.29795411303, 
    1760.03612032218, 
    1632.50565318022, 
    1613.38389819998, 
    1691.79874655368, 
    1450.65748871188, 
    1543.10237347936, 
    1586.55875170763, 
    1591.62384318944, 
    1389.0440088084, 
    1468.3059514524, 
    1402.12481161016, 
    1362.07719129383, 
    1234.71800419674, 
    1449.71098772245, 
    1249.36130939044, 
    1422.06447549034, 
    1242.45796069222, 
    1960.75750803998, 
    1764.43769455762, 
    1151.68574811023, 
    1351.94865847128, 
    1457.81826760554, 
    1584.64820561799, 
    1640.04120848664, 
    1735.31124281185, 
    1768.23630087453, 
    1918.99420702033, 
    1732.40993215134, 
    1760.0286585493, 
    1688.14273613463, 
    1772.07645690861, 
    1763.61924674239, 
    1740.11371863792, 
    1812.97517926928, 
    1770.18625833242, 
    1598.41125084341, 
    1697.48526766965, 
    1667.41316978565, 
    1867.52064941741, 
    1654.68895731847, 
    1749.52200898803, 
    1798.4252939017, 
    1959.43673495433, 
    1909.72233248543, 
    2012.91995125962, 
    2307.42546469999, 
    2246.58240490568, 
    2216.03158799454, 
    2384.55069244976, 
    2412.62701528326, 
    2425.99629235632, 
    2420.84859558385, 
    2369.14756348888, 
    2366.78761680882, 
    2288.37240773138, 
    2218.37698008831, 
    2106.87039240118, 
    2048.18741117175, 
    1975.04602125639, 
    1893.29571440982, 
    1875.78222008947, 
    1792.57159700643, 
    1728.25220098476, 
    1381.87824063449, 
    982.342213224737, 
    908.784102878628, 
    819.719442922024, 
    244.054277469676, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    660.559184950925, 
    861.480585150326, 
    952.208484885269, 
    1447.10605879639, 
    1308.91408856847, 
    716.256293605014, 
    971.751369673325, 
    1158.79792673457, 
    1644.10349590754, 
    1686.76262986256, 
    1714.29827181853, 
    2056.24812553746, 
    2023.84003788353, 
    1945.43741484042, 
    1904.65550526265, 
    1986.97310526439, 
    2069.80045993023, 
    2296.75559603706, 
    2361.08696199178, 
    2253.08289255152, 
    2177.49449531635, 
    2245.14275702109, 
    2220.12608538488, 
    2170.08379268521, 
    2222.92918621481, 
    2217.58501903799, 
    2029.58891248682, 
    1897.20472060718, 
    1734.52667580948, 
    1659.89280476319, 
    1797.12273328113, 
    1795.25718235392, 
    1800.35232187241, 
    1780.06375342241, 
    1683.4290284888, 
    1759.50644100346, 
    1700.39356854886, 
    1709.80577056811, 
    1681.35929519204, 
    1630.0462956031, 
    1597.16774557982, 
    1686.96831764089, 
    1681.13313705459, 
    1883.97422525228, 
    1812.11171094601, 
    1679.89131519127, 
    1702.79785523959, 
    1854.39702965775, 
    1789.1076377014, 
    1708.3712533354, 
    1694.36292733047, 
    1609.15569919914, 
    1734.09893662673, 
    1547.91528877628, 
    1578.85403636128, 
    1543.7671346329, 
    1601.09119913488, 
    1629.06920434711, 
    1707.7897229757, 
    1629.18815384621, 
    1545.31265586148, 
    1573.98012590638, 
    1623.83378705005, 
    1679.78104011357, 
    1985.1573077672, 
    1667.73868618063, 
    1519.69032903308, 
    1686.86183238307, 
    1905.26903153332, 
    1873.1010559186, 
    1920.51545650665, 
    1694.66798801755, 
    1781.58732274865, 
    1805.45575941234, 
    1806.86630439696, 
    1777.48646192251, 
    1757.23504073338, 
    1751.27944246501, 
    1883.71613186923, 
    1775.96533777887, 
    1902.8837477069, 
    1802.35231181663, 
    1706.30410691726, 
    1848.41711048511, 
    1892.91635169003, 
    2014.05035929846, 
    1782.98028656405, 
    1897.49078202871, 
    1999.60555831399, 
    2023.32478871845, 
    2097.3027270072, 
    2332.26545129929, 
    2367.59415111358, 
    2413.70448710389, 
    2410.24283481913, 
    2417.06737520843, 
    2461.05354704405, 
    2501.66299414621, 
    2469.91317977908, 
    2462.31469918468, 
    2468.31052209358, 
    2386.89880468336, 
    2318.60061298604, 
    2259.90804203801, 
    2210.05068743332, 
    2065.40322566918, 
    2031.16640979852, 
    1926.58336180935, 
    1826.163381953, 
    1625.81873998386, 
    1481.20321634407, 
    1339.75155581413, 
    1102.60683104939, 
    1158.54237470642, 
    1389.96510479282, 
    1187.86772879651, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    790.532533630118, 
    1142.2255784601, 
    1449.67075465401, 
    1238.51155033218, 
    1139.0055141576, 
    1024.83379513808, 
    1175.24219379398, 
    1668.54028984605, 
    1672.42389096355, 
    1939.34800192794, 
    2365.18930826027, 
    2267.45846119855, 
    1876.06036553607, 
    2104.69191589938, 
    1954.12663468235, 
    2168.58904475188, 
    2523.65055471728, 
    2517.68961954371, 
    2429.46682929821, 
    2330.42649511834, 
    2250.64372754255, 
    2175.21847357211, 
    2185.00199782241, 
    2307.67312121045, 
    2319.95211396285, 
    2214.73022969998, 
    1974.8559873512, 
    1843.92349148998, 
    1847.00965069785, 
    1866.65436916659, 
    1899.00183385758, 
    1934.51397880035, 
    1903.72868903923, 
    1874.83130031586, 
    1863.40663810918, 
    1874.84111480298, 
    1790.2591468137, 
    1737.87233849269, 
    1717.9312617861, 
    1733.98501739963, 
    1794.70920895763, 
    1909.35536318134, 
    1904.27357898915, 
    1907.93540634844, 
    1788.75465968574, 
    1834.95974409377, 
    2000.45577927186, 
    1823.79330982285, 
    2170.55569520606, 
    1939.67637071887, 
    1803.64292709572, 
    1709.22460120726, 
    1621.08819343867, 
    1556.93604829852, 
    1575.52625991672, 
    1556.71918525511, 
    1715.47589872597, 
    1707.88157264336, 
    1712.8511811001, 
    1730.946661247, 
    1708.56257437817, 
    1690.76180362664, 
    1501.58811605008, 
    1745.81784363705, 
    1834.16117629277, 
    1739.21749929495, 
    2047.99192342274, 
    2001.06034817582, 
    1867.4085955466, 
    1838.38437242156, 
    1820.1539526452, 
    1962.51911158748, 
    1955.9859423205, 
    1951.94397841592, 
    1928.2813538994, 
    2017.65715630614, 
    2023.25232717335, 
    1971.35295842716, 
    1898.29628480534, 
    1857.81600271708, 
    1764.26211902197, 
    1812.14191618266, 
    1955.03254403454, 
    2121.64399384805, 
    2095.27443789504, 
    2025.13971684348, 
    2129.45456674918, 
    2116.29618161887, 
    2042.02689630197, 
    2091.64117385712, 
    2404.84905948938, 
    2596.0284433605, 
    2570.26140693672, 
    2576.07892894188, 
    2564.38546561952, 
    2587.3629825448, 
    2580.46049304596, 
    2544.99273742557, 
    2548.01524238822, 
    2494.31176434904, 
    2502.24267927128, 
    2414.63239228703, 
    2328.51496044912, 
    2249.73105272833, 
    2204.11850292751, 
    2108.08618726448, 
    2045.39055074355, 
    1929.97720212149, 
    1812.48510241285, 
    1840.33861397521, 
    1551.32253947966, 
    1819.54715709852, 
    2088.48567881331, 
    1866.85137288318, 
    1077.1760452025, 
    618.468933835404, 
    0, 
    33.6671676961152, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    737.297507743053, 
    1166.11218347111, 
    965.843352351331, 
    1301.47201687022, 
    1347.00632426764, 
    1630.42469747785, 
    1718.27700332528, 
    1910.43728028846, 
    2145.82903040276, 
    2218.60656537468, 
    2332.42718520322, 
    2410.0469310155, 
    2376.10865092934, 
    2394.9342505707, 
    2562.56679827507, 
    2544.61333539728, 
    2485.60985110171, 
    2420.63522325147, 
    2300.93117133806, 
    2180.23370232901, 
    2123.97563812439, 
    2282.42703155846, 
    2226.4052707695, 
    2288.97118302989, 
    2167.63742246278, 
    2110.40159463074, 
    2083.74085603579, 
    2010.83941754061, 
    1993.48251521758, 
    2027.81114978226, 
    1972.85713098789, 
    1923.44175573379, 
    1989.5032648305, 
    1969.37198438824, 
    1939.0538636824, 
    1883.54458738152, 
    1867.90829969914, 
    1905.3831484163, 
    1906.59078716159, 
    1903.28864473211, 
    1942.1000371157, 
    2009.22289384313, 
    2041.96906400568, 
    1996.126402488, 
    1957.49588652875, 
    2027.85193760111, 
    2064.12512985206, 
    2022.33102110415, 
    1921.26266689531, 
    1966.43656152887, 
    1897.46900325832, 
    1757.30827833568, 
    1697.5268707927, 
    1783.69334712241, 
    1835.62383935641, 
    1828.93448431456, 
    1990.926338278, 
    1927.83614177161, 
    1848.85263065647, 
    1862.27391075399, 
    1741.5555597597, 
    1777.23037679517, 
    1991.3997595388, 
    2091.7669138536, 
    2013.77506239227, 
    2019.81281158762, 
    1927.59715160944, 
    1951.12639702272, 
    2030.19416031052, 
    2117.0907434016, 
    2104.04513372342, 
    2083.16585501033, 
    2063.85876057731, 
    2100.89346510582, 
    2162.80387665781, 
    2055.82196479149, 
    2034.97090860495, 
    1973.33360281065, 
    1924.3860051375, 
    1888.14298289992, 
    2146.04254167347, 
    2255.16777512831, 
    2222.27204175504, 
    2252.00970478663, 
    2298.15763496401, 
    2142.01083519591, 
    2097.91123425324, 
    2339.71785543593, 
    2552.112154841, 
    2710.40114971109, 
    2688.37394603828, 
    2641.36428335397, 
    2592.21825203639, 
    2712.90920793288, 
    2698.62131902462, 
    2638.8700253066, 
    2616.89609617967, 
    2595.40811832967, 
    2541.53977239636, 
    2548.19509122331, 
    2417.30825564475, 
    2305.23956530807, 
    2237.41759732423, 
    2175.46569994298, 
    2096.67520037235, 
    2064.25595355996, 
    2001.79630252193, 
    1996.89027563807, 
    1982.86810505494, 
    2033.64548026925, 
    1881.81136693974, 
    1323.72225997048, 
    1348.68718759024, 
    791.899332509333, 
    974.553953090462, 
    120.592766865798, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    887.185624307788, 
    717.335694104956, 
    815.777483306641, 
    790.09678014074, 
    1278.08387558325, 
    947.378115421115, 
    1659.05158190688, 
    1655.33422294007, 
    1779.32296182238, 
    2009.58445649364, 
    1890.48988536014, 
    1938.88512708986, 
    2080.01159358935, 
    2154.56197330008, 
    2467.53515261138, 
    2651.0992035478, 
    2525.54579579197, 
    2437.19289336498, 
    2532.37644133782, 
    2411.10971937226, 
    2218.48787312569, 
    2235.95196577607, 
    2200.27556408122, 
    2194.6360243447, 
    2287.32267267366, 
    2314.94285215604, 
    2389.21246901508, 
    2275.71545609417, 
    2197.20593465238, 
    2145.07397169966, 
    2169.94750291374, 
    2178.72723710786, 
    1990.42114472466, 
    2085.3624292233, 
    2052.23551296166, 
    2064.6439683473, 
    2056.02459477433, 
    2005.2116856954, 
    2130.45656957466, 
    2002.32279972393, 
    2042.19049941237, 
    2112.39862560037, 
    2153.47606556922, 
    2152.39632262141, 
    2111.85352741601, 
    2030.5497177504, 
    1986.00212544937, 
    2038.65124885786, 
    2163.71372462894, 
    2240.17314777171, 
    2199.38253459275, 
    2028.99702988837, 
    1987.96746017429, 
    1953.24777019139, 
    1997.16546798536, 
    1980.70558223825, 
    1990.28546113181, 
    2095.8959296983, 
    2083.24744435019, 
    2091.49371467334, 
    2084.25219488263, 
    2034.14074466371, 
    2127.359087844, 
    2245.73730026157, 
    2243.87216103279, 
    2144.99393499841, 
    2052.56925624129, 
    2037.07418581916, 
    2075.67284508492, 
    2165.50030780448, 
    2213.98971479923, 
    2222.31356452772, 
    2236.92184476298, 
    2239.74395606373, 
    2226.47586416178, 
    2255.88032098879, 
    2271.40752977752, 
    2290.57253385143, 
    2184.9383498017, 
    2161.10029784486, 
    2133.6734846371, 
    2204.26559067831, 
    2304.40189573109, 
    2331.14343004211, 
    2200.50627683839, 
    2418.72090102774, 
    2407.16423935268, 
    2531.41689953195, 
    2651.69684608385, 
    2637.21324359978, 
    2722.42744157731, 
    2661.85203465342, 
    2680.92848555687, 
    2763.20255556093, 
    2793.90241901752, 
    2793.50738334086, 
    2762.43600658997, 
    2731.85100673111, 
    2732.3353249275, 
    2635.18523555971, 
    2543.90131047617, 
    2459.86854335342, 
    2454.9893115235, 
    2343.81060491786, 
    2245.24184405234, 
    2168.04996375511, 
    2140.46360697357, 
    2121.40321625532, 
    2136.00222466519, 
    2139.88802732761, 
    1857.90311691284, 
    1479.00894423118, 
    1268.47335517597, 
    1242.47211676391, 
    965.536075668223, 
    801.957872229888, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    662.386429103705, 
    641.422517357733, 
    770.747062440825, 
    973.613652455038, 
    1262.50010783122, 
    1206.61692825157, 
    1884.06590420814, 
    1663.93043991162, 
    1582.44510971501, 
    1811.25753030679, 
    1697.96225895341, 
    1712.9448964095, 
    1745.06330959495, 
    2201.77499934107, 
    2564.00714721804, 
    2515.51256207223, 
    2415.26132324972, 
    2430.57421768451, 
    2688.87124462094, 
    2415.99141151242, 
    2254.22234133153, 
    2163.15541246185, 
    2077.41494881961, 
    2226.25401217141, 
    2325.75717359875, 
    2327.44778275471, 
    2325.92244645078, 
    2323.11635032119, 
    2282.08610710547, 
    2313.03481494796, 
    2294.75429918795, 
    2287.70411628209, 
    2243.87070661879, 
    2168.38470294976, 
    2188.08240325774, 
    2197.93094945106, 
    2179.30748788741, 
    2179.31536299173, 
    2179.3300440115, 
    2146.67214912388, 
    2139.67239532159, 
    2190.98782658397, 
    2146.9141533252, 
    2522.00485513609, 
    2349.14155300514, 
    2081.17739865522, 
    2196.80884116647, 
    2334.55704692318, 
    2178.20415533631, 
    2214.72022953405, 
    2263.69696337916, 
    2218.74206789939, 
    2211.1870265176, 
    2237.3800829219, 
    2175.43956372806, 
    2165.02017375383, 
    2275.54842113992, 
    2427.96439768279, 
    2335.56082126979, 
    1998.29658000643, 
    2124.80259617558, 
    2206.15711765238, 
    2436.60299986383, 
    2509.62675475646, 
    2356.41326301446, 
    2237.87138015578, 
    2139.27479109765, 
    2011.68870463523, 
    2232.89846234884, 
    2383.44076378087, 
    2409.18437927493, 
    2369.0542481693, 
    2347.51212521546, 
    2310.20289524677, 
    2344.53493599893, 
    2364.25771788938, 
    2455.31186590071, 
    2466.15265648223, 
    2396.16534754524, 
    2393.301013814, 
    2397.45874953668, 
    2336.34120591487, 
    2351.78832079663, 
    2308.61136541702, 
    2334.43392065362, 
    2531.09815080824, 
    2582.70144876488, 
    2647.89217322835, 
    2749.14968541467, 
    2775.0611700438, 
    2786.31487915746, 
    2768.73288988262, 
    2755.42260133212, 
    2859.19430059958, 
    2860.56302251554, 
    2839.34873069042, 
    2829.90915992467, 
    2798.54977800504, 
    2747.92859716802, 
    2674.49154212303, 
    2609.61262004543, 
    2592.84515442255, 
    2589.77526794286, 
    2435.953546774, 
    2333.15300955028, 
    2221.465869517, 
    2142.28333221886, 
    2182.13321300551, 
    2296.83372676283, 
    2200.92366886629, 
    1694.21235704391, 
    1490.65002774459, 
    1427.87514770316, 
    1273.21955608425, 
    787.269559759718, 
    640.134311749251, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    629.627942498031, 
    728.408672949556, 
    937.935469866244, 
    1153.84785264099, 
    1516.13384948979, 
    1650.38902495959, 
    1740.14319253338, 
    1607.17393311592, 
    1487.59556844023, 
    1531.65483823041, 
    1383.4773702233, 
    1643.06022360179, 
    1487.96881188944, 
    1807.46867381432, 
    2367.95985026039, 
    2243.9314802442, 
    2205.66661503128, 
    2320.01967052731, 
    2471.74323267294, 
    2309.83927674113, 
    2341.47581074756, 
    2084.77269606945, 
    2122.82211766077, 
    2405.5272777873, 
    2260.86713398585, 
    2376.75183813715, 
    2482.96089070395, 
    2311.00149249036, 
    2249.9268322121, 
    2287.51769671371, 
    2384.69449523054, 
    2419.59826979497, 
    2388.24972635775, 
    2323.74040325361, 
    2317.05231324784, 
    2324.38780674196, 
    2288.66733964252, 
    2298.91977600922, 
    2393.51315027663, 
    2314.01003278884, 
    2265.85337564115, 
    2239.06197382368, 
    2244.89653736121, 
    2313.76267750481, 
    2539.88052033249, 
    2279.41969857104, 
    2320.12364172701, 
    2396.83688148347, 
    2329.14027118456, 
    2256.29864686148, 
    2353.70499390195, 
    2470.39013920033, 
    2270.2275961058, 
    2282.09579093407, 
    2269.28466523777, 
    2298.86345500872, 
    2370.55724402836, 
    2295.36082606728, 
    2339.88638471585, 
    2116.22213080379, 
    2161.08174572999, 
    2279.06003570245, 
    2428.10606042455, 
    2492.21128837451, 
    2457.71132544282, 
    2340.52185166863, 
    2384.56186011638, 
    2394.35127695268, 
    2509.02507862449, 
    2625.31192997292, 
    2580.38843069184, 
    2599.69997306606, 
    2520.91229329493, 
    2487.55092641371, 
    2557.49137709841, 
    2559.72864588009, 
    2576.59439920662, 
    2654.73275279825, 
    2575.67325235242, 
    2553.66958246282, 
    2512.4710690509, 
    2463.3261061638, 
    2498.45133584928, 
    2479.48525041929, 
    2492.84616377519, 
    2542.83932031638, 
    2658.51661954326, 
    2734.3873438793, 
    2827.05012299376, 
    2872.93739417824, 
    2924.88437244553, 
    2904.14879016659, 
    2953.68430684025, 
    2951.84023353233, 
    2956.56739230941, 
    2923.95657012417, 
    2890.06002475573, 
    2854.33869412575, 
    2790.57423144547, 
    2727.66951237044, 
    2758.00680442852, 
    2731.29283354055, 
    2617.92177282513, 
    2522.95929831747, 
    2416.61608149697, 
    2310.62888415836, 
    2201.34527664983, 
    2145.72063335832, 
    2213.06833556915, 
    1932.79973266618, 
    1902.07332349789, 
    1505.60027130948, 
    1566.78294133048, 
    1098.48501964762, 
    692.383578733285, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1119.49663993816, 
    1002.73601703581, 
    779.241224640216, 
    668.576407524252, 
    1087.52380252794, 
    1173.22159546807, 
    1663.15181732254, 
    1411.50345792873, 
    1063.94567703759, 
    1393.87817838388, 
    1176.05243242902, 
    1084.03439232242, 
    1153.0377964281, 
    1862.23480296082, 
    2013.09956579372, 
    2039.73282720262, 
    2112.0715324914, 
    2342.90819543729, 
    2257.17950739219, 
    2245.43922198533, 
    2394.31428300677, 
    2122.89639727162, 
    2178.82837468551, 
    2001.9590058609, 
    2214.39419739402, 
    2507.51302623245, 
    2361.21367263285, 
    2245.24084452364, 
    2201.37774244215, 
    2371.19826205537, 
    2425.91810759278, 
    2460.09601676941, 
    2462.02644657278, 
    2409.92221982749, 
    2407.17875159858, 
    2381.07141414535, 
    2334.6716377413, 
    2312.87616356049, 
    2292.23651020992, 
    2360.1064212584, 
    2357.70783230881, 
    2333.17187743839, 
    2335.98806663061, 
    2476.37460938568, 
    2397.62798047113, 
    2155.45406043958, 
    2410.08196145723, 
    2493.56954464047, 
    2598.2446106588, 
    2557.64655578431, 
    2398.39052844126, 
    2549.40952896038, 
    2239.34662845677, 
    2271.12844182454, 
    2341.04536436666, 
    2365.34339503515, 
    2338.94434347879, 
    2262.2674016155, 
    2353.719852644, 
    2355.36292207306, 
    2357.4898290029, 
    2454.10011041452, 
    2549.86031538733, 
    2660.60323382801, 
    2638.47781166787, 
    2662.49396374263, 
    2638.79298694943, 
    2658.76278097906, 
    2656.49432534764, 
    2699.55008702468, 
    2646.3539417713, 
    2723.48422361785, 
    2706.38698507558, 
    2658.70189545989, 
    2665.95921179789, 
    2712.02133400729, 
    2722.56403602606, 
    2720.55306846024, 
    2595.66123900567, 
    2557.08958145664, 
    2516.52064470446, 
    2611.86700697071, 
    2653.34673219891, 
    2652.88205923887, 
    2638.17734939189, 
    2648.20451265798, 
    2713.3723424918, 
    2801.43126318389, 
    2915.34223546459, 
    2949.82220007791, 
    2964.85918972384, 
    2978.33424961805, 
    3010.0319794281, 
    2991.38301973542, 
    3014.97292334713, 
    2978.39965433555, 
    2964.1908615761, 
    2868.20861466503, 
    2828.77854821943, 
    2771.91263494545, 
    2759.93145555865, 
    2737.49586648148, 
    2678.75075929545, 
    2555.80179302224, 
    2419.86034443065, 
    2347.26057447656, 
    2234.85964187561, 
    2151.4418670621, 
    2330.46945733691, 
    1810.13920083028, 
    1917.10700491312, 
    1644.24162636257, 
    1394.93938643242, 
    1116.78214349638, 
    896.547733284246, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    727.505004349355, 
    904.671174478137, 
    874.679769172174, 
    897.184994383386, 
    951.20538594615, 
    545.043635990281, 
    1212.45928004791, 
    1177.87678863847, 
    694.698372503499, 
    1143.95990642697, 
    1520.85477436589, 
    1197.11318862804, 
    1146.99567514253, 
    1489.1297215687, 
    1675.32947856249, 
    1937.58460128317, 
    2171.68694841519, 
    2338.91835692776, 
    2099.73256166215, 
    2137.78281293361, 
    1963.96368982121, 
    1981.45919646485, 
    1982.8145331836, 
    2056.03283415635, 
    2328.07402895984, 
    2464.28886459416, 
    2397.17782537155, 
    2283.53895634455, 
    2272.53534756828, 
    2371.65865706294, 
    2456.44635008781, 
    2445.81436197596, 
    2520.53481875586, 
    2517.70122956751, 
    2441.44980649121, 
    2425.09604545072, 
    2403.8744274698, 
    2377.89226714416, 
    2402.33676415131, 
    2434.82097034468, 
    2434.12882281005, 
    2430.26813123325, 
    2464.4730096877, 
    2527.8099444757, 
    2430.69157568291, 
    2445.10282909996, 
    2422.37670025776, 
    2478.51561950104, 
    2663.73093969556, 
    2468.15906725791, 
    2412.05200123776, 
    2484.26861422007, 
    2423.40373455004, 
    2492.14258495829, 
    2622.30316082949, 
    2669.11468795173, 
    2491.91138047089, 
    2449.64552645529, 
    2478.35441712193, 
    2591.36722711236, 
    2500.50543711421, 
    2659.54198392034, 
    2666.03291295119, 
    2720.52064494341, 
    2777.72813398236, 
    2866.62062148838, 
    2808.82919667903, 
    2814.69194442123, 
    2731.70302387886, 
    2781.73643346404, 
    2756.85522507487, 
    2833.68611884728, 
    2866.48355183367, 
    2784.7590347183, 
    2745.42926696067, 
    2843.97423264555, 
    2785.48727647106, 
    2695.97361018772, 
    2685.03665941543, 
    2702.10857574397, 
    2744.47582450997, 
    2868.51745727781, 
    2882.27994728571, 
    2880.78293555913, 
    2809.38390160285, 
    2781.76483592113, 
    2845.4901704517, 
    2897.83631369981, 
    2947.76418944776, 
    3002.77122906871, 
    3071.57614710239, 
    3072.14364331474, 
    3092.27584098042, 
    3094.99694549037, 
    3090.30893753693, 
    3037.57980944386, 
    3052.06148789377, 
    2962.56832667665, 
    2892.08280766034, 
    2850.96586425939, 
    2795.27921701675, 
    2755.22150276348, 
    2652.57487412901, 
    2548.95493739192, 
    2476.93941576295, 
    2341.44092024764, 
    2213.10773623546, 
    2107.64518554516, 
    2220.5326326868, 
    2065.55096725339, 
    1948.38495411569, 
    1820.28356164853, 
    1704.39827815557, 
    1424.64421902247, 
    971.958631869894, 
    1208.90304403136, 
    28.7797698470213, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1035.19782806302, 
    656.182910310492, 
    603.074539303963, 
    1150.64562093465, 
    772.453966261729, 
    792.063088489252, 
    726.523763127032, 
    1159.35106024486, 
    953.676106557678, 
    1116.79181174526, 
    1167.86537736513, 
    868.632155804553, 
    1143.05559162597, 
    1334.21511037319, 
    1428.96325718658, 
    1559.99702473827, 
    1770.15454914251, 
    1809.17949865366, 
    1806.97100703108, 
    1846.31948463541, 
    1829.68565735917, 
    1864.97496898282, 
    2099.3857104693, 
    2253.34467676221, 
    2074.38292166957, 
    2264.80866009664, 
    2429.02675433753, 
    2265.78726467337, 
    2208.74651507026, 
    2274.70800497529, 
    2474.79803246718, 
    2571.49305831098, 
    2562.49008203004, 
    2554.3893338743, 
    2538.14446975555, 
    2554.42166185988, 
    2475.68055125327, 
    2441.62736165917, 
    2514.26016767262, 
    2601.88172920046, 
    2554.91787570037, 
    2511.45751051725, 
    2442.36345590601, 
    2558.92337638821, 
    2548.72331844673, 
    2582.06009069907, 
    2538.15793850656, 
    2590.9997444348, 
    2679.21931567766, 
    2510.47383769524, 
    2654.77891727642, 
    2629.11728698716, 
    2564.48233051906, 
    2682.88205346524, 
    2826.88868747031, 
    2866.77049740825, 
    2710.89515865194, 
    2664.55909358262, 
    2632.74733005326, 
    2581.23848415494, 
    2598.59631066856, 
    2706.34809187355, 
    2814.29683193979, 
    2898.57391529228, 
    2931.20955529084, 
    2944.75930888944, 
    2948.31626495818, 
    2949.85239069157, 
    2931.9095740068, 
    2900.65561330752, 
    2851.83841672828, 
    2938.14856157442, 
    2946.27494937794, 
    2924.50986256534, 
    2913.85772504037, 
    2972.77264321094, 
    2818.34790633434, 
    2750.43929891792, 
    2796.87863362366, 
    2897.0013714024, 
    2970.0019576059, 
    2918.3898902969, 
    2992.44798690137, 
    3078.43417275973, 
    2873.20858358368, 
    2916.01910458079, 
    3042.3633568138, 
    2933.30498015562, 
    3033.39136784286, 
    3110.70450894176, 
    3140.11534712148, 
    3142.10986201518, 
    3225.76803755075, 
    3119.74296712642, 
    3113.77393344981, 
    3116.7957481881, 
    3077.48217376901, 
    3047.26462996103, 
    2956.8865621899, 
    2868.95223484236, 
    2795.66446793879, 
    2730.85329783461, 
    2669.29271008884, 
    2520.76701648942, 
    2440.18434949613, 
    2313.48466977391, 
    2148.14825801516, 
    2184.75832379603, 
    2313.75309313853, 
    1923.71552448481, 
    1798.11048615883, 
    1502.8812506395, 
    1366.90004691158, 
    1130.00201780487, 
    839.763434696596, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1073.21328058247, 
    827.189671260353, 
    627.754485112721, 
    954.267922783981, 
    760.572351250554, 
    808.073127521993, 
    854.042488174713, 
    1518.14946384723, 
    1517.27000573263, 
    961.921297684294, 
    1009.30462881903, 
    580.584461139018, 
    815.907415065206, 
    1243.89974066757, 
    1084.14138846346, 
    1478.20793775583, 
    1502.22118153451, 
    1315.77932121287, 
    1385.49421079243, 
    1791.85392533702, 
    1589.06926658664, 
    1810.62444960813, 
    1872.06239972762, 
    1793.34529150286, 
    2090.95736248898, 
    2233.83070016614, 
    2126.6760148436, 
    2023.07956053374, 
    2367.89489691783, 
    2540.31962617766, 
    2626.73328011987, 
    2648.55410982196, 
    2614.13054520046, 
    2565.65777005805, 
    2532.41448777352, 
    2532.12830621571, 
    2507.55964230423, 
    2576.42632571809, 
    2585.83963075501, 
    2613.13374846063, 
    2652.53749533999, 
    2747.8572003864, 
    2649.7926153369, 
    2736.78568289337, 
    2689.58865490713, 
    2664.92718993203, 
    2759.73762105771, 
    2738.10556901204, 
    2581.16391069362, 
    2693.0773888993, 
    2752.76135341604, 
    2577.74116397618, 
    2658.32884496587, 
    2803.38225796977, 
    2815.81428306282, 
    2787.52926431339, 
    2786.8675067814, 
    2766.52053483064, 
    2754.77071974016, 
    2731.7987414207, 
    2786.45093003976, 
    2956.38083738407, 
    3064.2113748493, 
    3062.17645735337, 
    3039.48415713327, 
    3081.96783338611, 
    3112.20134085002, 
    3081.36185260159, 
    3017.44444590535, 
    3052.67325342805, 
    3061.19689588402, 
    3047.79489028956, 
    3056.82164806853, 
    3006.87699390238, 
    3051.34865920328, 
    3024.43392029816, 
    2939.20880636871, 
    2957.49563021966, 
    2996.44912186695, 
    2954.20181287236, 
    2980.12853964125, 
    3024.26905328373, 
    3050.11842933525, 
    2990.4327052594, 
    3083.20064697531, 
    3240.13940903339, 
    2997.49544544969, 
    3092.6182748023, 
    3207.89152289296, 
    3084.03095842606, 
    3171.63001098038, 
    3181.22466205916, 
    3165.66934989247, 
    3143.92520296336, 
    3078.0222898714, 
    3083.59514696085, 
    3092.3686070495, 
    3090.46687078572, 
    2900.47316244518, 
    2772.59059831143, 
    2763.59353119222, 
    2678.86981904044, 
    2705.75724363447, 
    2751.3703290157, 
    2639.48622788751, 
    2477.84554813384, 
    2444.52897991152, 
    2121.74581901382, 
    1871.150713626, 
    1704.89683971706, 
    1586.59517185125, 
    1419.52462445669, 
    1169.97123293237, 
    876.539419602374, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    869.376638163946, 
    717.12109547268, 
    820.019300021224, 
    922.380751522692, 
    1083.18647449186, 
    885.465687297499, 
    1390.80004069391, 
    1295.33872349432, 
    680.487607497193, 
    741.657133928953, 
    1271.07571298996, 
    737.140329762793, 
    789.603294959563, 
    1076.70869863229, 
    1369.82012243596, 
    1098.48172007299, 
    1306.96072902564, 
    1619.45865633114, 
    1550.27577709473, 
    1555.11161618757, 
    1565.31772251696, 
    1959.13633643206, 
    1954.21048455701, 
    1938.35047187012, 
    2011.70569954838, 
    2102.71368200594, 
    2214.25499849466, 
    2370.46777078713, 
    2577.60262282194, 
    2670.08609970997, 
    2482.80038616165, 
    2593.67677560997, 
    2689.97406615418, 
    2624.51126140651, 
    2629.47851551501, 
    2601.79338270088, 
    2564.12034611977, 
    2648.84782264908, 
    2729.99607954561, 
    2803.34613198456, 
    2803.93826643791, 
    2710.04021081018, 
    2664.49013046835, 
    2693.73647509115, 
    2791.62390849607, 
    2755.94734699729, 
    2728.5296087638, 
    2743.00417969807, 
    2736.67411210435, 
    2718.75439102345, 
    2700.9171006051, 
    2773.7879677441, 
    2814.13191873754, 
    2841.69885010349, 
    2907.63218747532, 
    2876.10608057209, 
    2860.77622752043, 
    2924.39837777887, 
    2990.98596443408, 
    3096.77391457088, 
    3192.46996026256, 
    3197.06975863445, 
    3142.24740229197, 
    3165.5963506841, 
    3295.34477149595, 
    3250.29143179961, 
    3189.80924298273, 
    3206.50035828736, 
    3158.78939727319, 
    3151.72216445155, 
    3126.64324935101, 
    3117.88972100375, 
    3128.53435945666, 
    3137.77340980256, 
    3100.06363918702, 
    3067.49709958326, 
    3053.48247272662, 
    3066.97496324319, 
    3110.83606889286, 
    3125.80248948241, 
    3157.5495068465, 
    3185.30746162974, 
    3213.56176451337, 
    3191.76175416909, 
    3203.98325010477, 
    3161.02134546482, 
    3203.55110528038, 
    3163.00711346703, 
    3268.05485006756, 
    3167.13193123644, 
    3206.70657578718, 
    3181.79556495263, 
    3071.70888625255, 
    3094.9544813413, 
    3038.4458754116, 
    3019.16772193565, 
    2933.7463117585, 
    2850.56708404523, 
    2795.83310764379, 
    2742.31603044935, 
    2675.01537286812, 
    2531.57205886945, 
    2336.3466687865, 
    2410.91720888762, 
    2252.92405832775, 
    2220.12349900181, 
    1996.06085212991, 
    1713.62251545243, 
    1685.67268964479, 
    1878.6139899209, 
    2037.60326115885, 
    1802.0807451338, 
    1299.24280505206, 
    0, 
    87.40478515625, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1122.65130476611, 
    663.80313214819, 
    1146.07728697404, 
    1280.9828447711, 
    722.324553703151, 
    819.70531100482, 
    739.697376523492, 
    892.389975507114, 
    1318.99023772806, 
    1290.36408680629, 
    1442.89289043944, 
    1388.33984929919, 
    1735.41189940887, 
    1443.93522877642, 
    1394.40193243889, 
    2008.94183517103, 
    1808.15155986162, 
    1968.68355567783, 
    2028.14495428843, 
    2199.96284399514, 
    2333.19855271596, 
    2383.13689565519, 
    2480.39140318641, 
    2519.78463176736, 
    2397.39229383993, 
    2548.2615283023, 
    2575.69286295523, 
    2654.02231469184, 
    2727.20025409285, 
    2635.12848945517, 
    2660.34443021412, 
    2743.32330049049, 
    2764.42986478652, 
    2836.31809545663, 
    2908.56935113169, 
    2789.17315533359, 
    2788.0835502567, 
    2799.65275915136, 
    2782.42087098986, 
    2744.9386745183, 
    2728.85227342715, 
    2732.03403597109, 
    2774.43801830505, 
    2760.47712176017, 
    2784.43788144954, 
    2857.66184110064, 
    2878.86059036612, 
    2917.29480762724, 
    2930.76073297842, 
    2916.60612475403, 
    2952.7746053199, 
    3024.84640287623, 
    3097.47288291773, 
    3205.82549848867, 
    3293.44706745513, 
    3294.60550106592, 
    3273.78510127962, 
    3314.8409638837, 
    3392.19600366792, 
    3409.74747895073, 
    3379.48129919276, 
    3353.94514324644, 
    3358.05030650265, 
    3301.0694200388, 
    3286.41711156885, 
    3249.46414336609, 
    3218.52231221404, 
    3206.65148485534, 
    3172.320210594, 
    3170.49391279485, 
    3154.30032209706, 
    3164.77443334259, 
    3271.85714580936, 
    3306.62701448909, 
    3334.52862653394, 
    3333.46871976079, 
    3314.4401494657, 
    3333.82096287417, 
    3251.51993515432, 
    3231.62178545735, 
    3271.67683615937, 
    3343.4910220974, 
    3146.63247298523, 
    3147.53505068789, 
    3193.28748649046, 
    3180.47284133138, 
    3146.18715401772, 
    3117.58860055856, 
    3033.16694621621, 
    3018.62836573001, 
    3007.5147041432, 
    2957.00437773978, 
    2860.31623404838, 
    2835.49983351338, 
    2656.58621707013, 
    2543.17372415512, 
    2467.29133942313, 
    2435.07574265075, 
    2319.65717301391, 
    2254.23927622274, 
    2116.12309330222, 
    1779.64219811454, 
    1692.94350129129, 
    1814.7282668264, 
    1326.54441400538, 
    964.0066674273, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    521.146494421645, 
    1084.81113100083, 
    1278.448059424, 
    821.193770942824, 
    1188.45810658985, 
    960.493219754431, 
    1394.05818150753, 
    1236.50449378051, 
    1234.44953164581, 
    1248.51732143839, 
    923.531378942907, 
    1675.55429477147, 
    1669.62673981189, 
    1801.0819207397, 
    1888.59509974907, 
    1978.75529279575, 
    2102.22185882964, 
    2145.16198605604, 
    2241.58605895672, 
    2480.03575864186, 
    2570.17379729484, 
    2578.48265969524, 
    2631.58102680724, 
    2696.98794246245, 
    2752.3413861434, 
    2672.28216513632, 
    2814.54465305611, 
    2709.58858526938, 
    2747.07200341507, 
    2752.7405100498, 
    2769.74585511065, 
    2928.50928341377, 
    2880.53095211703, 
    2956.619517968, 
    2940.03567675522, 
    2852.81086013523, 
    2808.39910608923, 
    2769.19661212867, 
    2759.22414123138, 
    2777.36953311135, 
    2804.92874641586, 
    2880.02428173217, 
    2935.07894653229, 
    2929.61673554306, 
    3040.96902527739, 
    3060.44170143091, 
    3036.1920055531, 
    3019.74822698278, 
    3102.23253960351, 
    3178.02177256412, 
    3261.62436063643, 
    3304.71384597898, 
    3345.07810651893, 
    3449.74270301945, 
    3243.06769257167, 
    3343.87989415654, 
    3389.31107068312, 
    3416.39688130093, 
    3503.2823534531, 
    3603.67134950496, 
    3540.62469258734, 
    3444.28116805547, 
    3329.06473999481, 
    3302.2474947077, 
    3298.30322390255, 
    3273.55462471478, 
    3286.26466329654, 
    3302.33743072088, 
    3355.10601944889, 
    3384.12468947812, 
    3361.93826150724, 
    3342.79597761551, 
    3334.68751332231, 
    3360.05846101095, 
    3412.54098061385, 
    3323.79227776008, 
    3362.66146642705, 
    3197.00647775209, 
    3167.59779965614, 
    3169.44576917276, 
    3173.89330383159, 
    3167.7411114936, 
    3312.62919941124, 
    3139.85212837009, 
    3073.16390359375, 
    3017.77883296221, 
    3019.77263707818, 
    3042.42045765158, 
    2985.95721620768, 
    2888.48885720432, 
    2802.32358707493, 
    2687.81637243073, 
    2562.40137216662, 
    2536.75939022737, 
    2486.91731364726, 
    2378.91920957026, 
    2125.89137680634, 
    1881.81412910047, 
    1857.02933869678, 
    1728.99005489085, 
    1447.17629082506, 
    1393.49494640035, 
    1117.45422264352, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    894.72323907076, 
    1055.98527918246, 
    722.303926127211, 
    1282.6694252335, 
    1108.76669726403, 
    910.501739958409, 
    1782.94190847712, 
    848.776688438769, 
    799.668795869934, 
    1018.15382861958, 
    1378.45833334364, 
    1447.68092267813, 
    1455.73846125285, 
    1746.55215572054, 
    1858.42255220106, 
    1986.91310753124, 
    2037.61581381818, 
    2253.9507005586, 
    2337.57325172521, 
    2379.72089139976, 
    2396.59589717098, 
    2508.07413245663, 
    2609.65358745117, 
    2729.18962417874, 
    2849.48340647192, 
    2846.50562929689, 
    2936.08006612831, 
    2923.76643543593, 
    2909.12644627209, 
    2849.25113478295, 
    2687.01918664316, 
    2922.96577508395, 
    2846.66769067264, 
    2869.83385519301, 
    2962.18580189876, 
    2926.62564575948, 
    2891.3551150361, 
    2821.42153970825, 
    2841.08408722288, 
    2940.64305325978, 
    2952.0393966152, 
    2910.59396960804, 
    3055.69046385249, 
    3082.17041214884, 
    3172.69794405602, 
    3103.2086629748, 
    3077.07183436561, 
    3124.30648206248, 
    3130.16316873604, 
    3254.1471518841, 
    3322.17445317303, 
    3373.05077850139, 
    3424.03258938975, 
    3365.16116158886, 
    3411.42476876537, 
    3424.47260358877, 
    3450.72176378785, 
    3382.27911631119, 
    3398.57108972058, 
    3422.50234697877, 
    3438.29976826418, 
    3472.61951366842, 
    3381.06763891829, 
    3400.95327003296, 
    3427.52637508519, 
    3440.93193062861, 
    3509.16979784628, 
    3517.36800296453, 
    3412.8869808536, 
    3407.460128797, 
    3415.17381833471, 
    3411.0907718337, 
    3425.66744402146, 
    3377.55248371764, 
    3320.44959511765, 
    3312.11684602792, 
    3311.66542165453, 
    3286.77987665192, 
    3273.21180647387, 
    3201.44973725416, 
    3213.5143474243, 
    3188.10508242051, 
    3222.65422085412, 
    3099.97855526822, 
    3012.65203757814, 
    2982.41902401056, 
    2978.62989809012, 
    2965.17038189746, 
    2935.75392202845, 
    2909.8351752748, 
    2809.35671372411, 
    2684.47687420424, 
    2554.87425113951, 
    2456.93010275166, 
    2388.05067348758, 
    2347.3072375515, 
    2151.66016299903, 
    1961.47544591606, 
    1864.46651058164, 
    1600.5359704295, 
    1368.93097126829, 
    1183.23008853219, 
    1038.71886474361, 
    775.2176386971, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    981.716865960341, 
    668.079638245746, 
    538.495748124623, 
    526.748658270962, 
    1309.05293735964, 
    1446.77265219078, 
    709.977643054881, 
    682.502811588632, 
    1032.61139234851, 
    1394.05412059069, 
    1348.72927030695, 
    1343.43349844513, 
    1720.00278162845, 
    1776.8218378123, 
    1892.41062961423, 
    2054.52736249379, 
    2192.94178496444, 
    2183.52570775386, 
    2198.51272306007, 
    2298.74649950389, 
    2492.43291626461, 
    2566.81997866317, 
    2738.66522398197, 
    2763.76173698577, 
    2756.45442324213, 
    2866.62254576127, 
    2929.16148596931, 
    2904.87989030132, 
    2938.63808184074, 
    2994.96254765806, 
    3008.27025337293, 
    2805.19486708169, 
    2920.97889859838, 
    3111.06733028533, 
    2978.57460387396, 
    2920.22160268948, 
    2816.57799245666, 
    2946.7914276883, 
    3082.87404194695, 
    3018.65970172881, 
    2971.86608758135, 
    3135.63719593431, 
    3219.54058795198, 
    3203.49469723068, 
    3142.16569049586, 
    3139.3818658568, 
    3216.12983963101, 
    3227.57388962011, 
    3329.89714150935, 
    3411.07539630552, 
    3452.60759930572, 
    3450.4199965215, 
    3373.71413841428, 
    3491.47642133694, 
    3482.60813918173, 
    3417.62093109961, 
    3409.67917806594, 
    3419.18243886843, 
    3416.53193064848, 
    3464.88837617257, 
    3492.03948812288, 
    3493.88752923589, 
    3514.33145430995, 
    3484.48410236321, 
    3483.36824108115, 
    3461.90547423831, 
    3457.43808066932, 
    3430.45059895606, 
    3443.65361919222, 
    3444.33754953192, 
    3419.29601808706, 
    3420.17407951093, 
    3371.54317960569, 
    3345.45443350266, 
    3342.41866176457, 
    3348.14380278708, 
    3324.41572252313, 
    3286.83971988472, 
    3239.14065643808, 
    3204.16887492317, 
    3165.48538355017, 
    3154.07563247963, 
    3050.01700768466, 
    3039.14377047641, 
    3011.22208591193, 
    3001.4227424065, 
    2986.98824475419, 
    2946.76197805068, 
    2888.73865292997, 
    2820.20980561644, 
    2726.96360913777, 
    2522.3844813072, 
    2459.59924021265, 
    2485.30109517618, 
    2377.10926097545, 
    2290.00137839033, 
    2087.76458030398, 
    1830.14787606643, 
    1710.30584403347, 
    1634.94867530761, 
    1389.05432921714, 
    1557.76294436234, 
    1428.24190854989, 
    573.319258823313, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    955.057589740113, 
    1180.42946784405, 
    976.556032749735, 
    1221.00972066573, 
    963.392676049458, 
    692.413844198804, 
    1052.05198071235, 
    0, 
    1341.73247890814, 
    1142.42314314375, 
    1392.66254287919, 
    1586.07155565224, 
    1741.221267522, 
    1982.27016874712, 
    2021.42452693492, 
    2060.48872627934, 
    2244.45592833084, 
    2369.31561721411, 
    2493.00332778453, 
    2661.8832354424, 
    2753.66082651508, 
    2707.8736028669, 
    2687.77258973359, 
    2804.28117546998, 
    2980.52453205151, 
    2969.23550031454, 
    3065.42628961986, 
    3103.26250684294, 
    2999.76763696807, 
    2868.00048036938, 
    2969.61894377815, 
    3099.23034501703, 
    3041.38805362836, 
    2962.35917798744, 
    2954.83040499103, 
    2997.28225690515, 
    3085.28847352626, 
    3073.41157497528, 
    3034.16382577816, 
    3055.61141969096, 
    3133.09822968204, 
    3254.12455002496, 
    3220.85424089971, 
    3199.6972854897, 
    3244.70865528806, 
    3343.33004713029, 
    3406.90243753947, 
    3472.64567308615, 
    3480.53998955634, 
    3465.40634058092, 
    3435.2992939711, 
    3390.60161694133, 
    3385.56420643679, 
    3404.89783218542, 
    3434.97322806163, 
    3454.61353642028, 
    3494.29479094179, 
    3553.1114551437, 
    3579.16911480145, 
    3564.30785263478, 
    3569.0401850546, 
    3520.79934858858, 
    3492.62331422251, 
    3490.24691612515, 
    3486.82521584755, 
    3459.37667646811, 
    3442.53553815181, 
    3435.39591164094, 
    3371.61671369449, 
    3393.01669607157, 
    3366.23757533395, 
    3346.14599664267, 
    3345.87632261401, 
    3342.2143536084, 
    3328.1754782017, 
    3299.25405743095, 
    3245.55004536909, 
    3180.44516563156, 
    3161.39767119735, 
    3198.41327142825, 
    3051.96380824888, 
    3035.34962986684, 
    3000.71520448501, 
    2990.94996251449, 
    3008.89752219968, 
    2914.12647552169, 
    2861.78763021924, 
    2821.23523976992, 
    2769.3408510221, 
    2641.80804732188, 
    2552.89023823923, 
    2477.23953820105, 
    2326.85049309692, 
    2284.52324429968, 
    2058.06918806269, 
    1890.72434405558, 
    1826.34102857167, 
    1607.96062862421, 
    1492.70806742859, 
    1171.52789957251, 
    1015.678403184, 
    801.602790263618, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    731.427705086704, 
    0, 
    0, 
    939.994167944581, 
    860.815268565159, 
    822.319990276052, 
    1150.79131795955, 
    1492.77956713196, 
    1530.45263578416, 
    1676.76184826802, 
    1851.00979395973, 
    2176.80562640186, 
    2292.71423921056, 
    2415.29581244348, 
    2569.89186209999, 
    2592.92555049913, 
    2692.53703727794, 
    2637.02790568371, 
    2562.2166944477, 
    2774.27631526209, 
    3000.62289906448, 
    3079.50944928955, 
    3094.46932968781, 
    3136.92600805423, 
    3057.66916440832, 
    3011.23281475502, 
    2984.65656657536, 
    2937.67420758133, 
    3006.7436500431, 
    3088.70175002901, 
    3239.82375098894, 
    3139.23388581019, 
    3208.97779299759, 
    3199.64929633346, 
    3112.14410016162, 
    3085.30454343803, 
    3218.64169171725, 
    3305.28872614088, 
    3216.75277780838, 
    3278.89371205265, 
    3334.04176989452, 
    3376.5533653048, 
    3432.30354204396, 
    3499.38207737303, 
    3476.45418749226, 
    3450.9122566685, 
    3320.8938313448, 
    3373.00726794127, 
    3350.93709822686, 
    3377.93892260549, 
    3526.98225950926, 
    3421.00034656537, 
    3552.77145929672, 
    3592.16879925123, 
    3612.78177775882, 
    3613.57415099899, 
    3593.38731986054, 
    3550.58907386146, 
    3486.04081350988, 
    3430.02281509039, 
    3465.27469364782, 
    3448.10815584148, 
    3450.91180953678, 
    3427.10003273568, 
    3362.89746554575, 
    3388.31276444348, 
    3387.11713863335, 
    3351.04617956734, 
    3334.36023382073, 
    3335.81533755051, 
    3293.12214646518, 
    3247.26024891106, 
    3228.19411450937, 
    3157.39383011735, 
    3119.26022009157, 
    3132.78765988481, 
    3062.43731301051, 
    3016.37586904227, 
    2913.40724401211, 
    2865.45579340441, 
    2825.91917437811, 
    2847.25516530319, 
    2828.16912291487, 
    2767.88572573589, 
    2756.61478068316, 
    2726.59429623648, 
    2644.14074565012, 
    2554.00812101513, 
    2451.62195225961, 
    2239.25533879573, 
    2072.39212992039, 
    1823.12204671271, 
    1693.47784403563, 
    1574.0048530991, 
    1195.33346215366, 
    945.530445754935, 
    871.953732227326, 
    1194.41120442033, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1160.35622692371, 
    993.808812459065, 
    1455.69999191619, 
    1346.29093686112, 
    1432.04833329906, 
    1632.31286680313, 
    1794.74426965426, 
    1842.24864863655, 
    2095.81142050594, 
    2313.14432582206, 
    2428.95798752903, 
    2346.52436875851, 
    2550.60128400705, 
    2672.80717251149, 
    2812.54216767278, 
    2885.39313096251, 
    3019.20509896439, 
    3192.74284723368, 
    3190.39018686354, 
    3172.15967750875, 
    3096.62868752562, 
    3011.05559084622, 
    3006.83863165679, 
    3114.10399111109, 
    3079.34830133077, 
    3095.07529328025, 
    3288.38379985376, 
    3216.35168391199, 
    3201.39530232712, 
    3237.23441771849, 
    3244.8850868369, 
    3315.34894924166, 
    3325.30372102041, 
    3294.82155715195, 
    3153.00425701068, 
    3299.02770839673, 
    3372.69953306862, 
    3413.51117265397, 
    3473.1488364462, 
    3492.52853716869, 
    3495.22341623245, 
    3466.18801039034, 
    3406.86800247661, 
    3411.65247312959, 
    3343.41216146098, 
    3350.40709768796, 
    3468.82381606208, 
    3478.36223902086, 
    3534.35266895883, 
    3640.38380100704, 
    3646.4698068053, 
    3627.40387083025, 
    3583.92550496839, 
    3513.44887947684, 
    3488.77206370078, 
    3434.19870884564, 
    3459.54530130171, 
    3426.23359162834, 
    3445.01690749695, 
    3392.59660896749, 
    3346.67471408873, 
    3344.07930689388, 
    3322.35406496536, 
    3313.65650604881, 
    3252.55764977464, 
    3273.27405194298, 
    3237.67007262085, 
    3210.55316490983, 
    3192.22309309784, 
    3110.48456733828, 
    3096.76965673831, 
    3180.02569697331, 
    3125.79887106553, 
    3027.65301169426, 
    2848.72861591255, 
    2952.09926668907, 
    2796.67890239312, 
    2817.8888104392, 
    2788.76194058417, 
    2763.15601453271, 
    2744.51114958297, 
    2705.76457714828, 
    2620.29668392147, 
    2585.5607952693, 
    2440.66948661636, 
    2151.65127854234, 
    2058.37827752701, 
    1949.0542584918, 
    1742.98962743838, 
    1614.3867943789, 
    1405.51943623923, 
    1083.78506192422, 
    899.784743550859, 
    922.617792600523, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    954.683641108239, 
    0, 
    1039.17582845712, 
    1131.31843974471, 
    1407.25235814771, 
    1723.33361350496, 
    1941.71280440377, 
    2095.34389788116, 
    2209.40643876001, 
    2269.8853712876, 
    2389.78204915678, 
    2364.99342774719, 
    2718.77273922036, 
    2924.53029675378, 
    2953.34981224406, 
    2901.37119469147, 
    2968.34275570936, 
    3025.31288000053, 
    3091.18362962138, 
    3102.68550463153, 
    3127.05978307854, 
    3202.68560461298, 
    3157.78748455777, 
    3153.89502212279, 
    3208.58460052377, 
    3281.78415416589, 
    3191.76490745828, 
    3203.07937992059, 
    3248.60768190952, 
    3300.44393708283, 
    3346.60047997932, 
    3366.16911180124, 
    3305.61998347098, 
    3232.10354687168, 
    3256.85413083315, 
    3342.75938929933, 
    3522.51401879266, 
    3578.4443439089, 
    3518.64511630872, 
    3466.09508016024, 
    3453.55316536558, 
    3398.85142566936, 
    3450.94698434399, 
    3467.96279494385, 
    3379.0805760654, 
    3452.69482894179, 
    3525.34016477572, 
    3560.88494088008, 
    3634.44090325753, 
    3700.09063063357, 
    3604.37234748988, 
    3558.48825629132, 
    3502.46655168771, 
    3490.74055276881, 
    3429.38902358203, 
    3461.97160375773, 
    3442.25098100971, 
    3390.4775032791, 
    3337.11063406355, 
    3295.9688872058, 
    3262.35558611503, 
    3247.62364540429, 
    3204.35910003854, 
    3115.51929736858, 
    3101.72202187116, 
    3134.53014321468, 
    3158.94351989298, 
    3149.8334190697, 
    3081.93549508663, 
    3001.98587044135, 
    3018.89819836181, 
    3055.4950428656, 
    2949.34413327842, 
    2764.86089522222, 
    2892.61795431937, 
    2765.37429400867, 
    2763.24135146403, 
    2795.23546949051, 
    2672.85674222157, 
    2652.82934788145, 
    2617.59138139925, 
    2537.30668232641, 
    2507.74341858158, 
    2478.00301833678, 
    2366.96695908467, 
    2212.35829350285, 
    2062.92081320785, 
    1798.3056422767, 
    1623.2938793023, 
    1588.58784785508, 
    1270.36298868937, 
    1045.31940593815, 
    833.500799615095, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1021.88342050919, 
    1027.53336867074, 
    853.938875898934, 
    1146.40296914558, 
    1496.80741683077, 
    1909.99413317057, 
    2105.15840402626, 
    2114.331500504, 
    2122.5527627818, 
    2131.34804647259, 
    2455.39956326281, 
    2676.55604459041, 
    2897.07356568634, 
    2953.00866167769, 
    2967.80948136278, 
    2879.19149302452, 
    2857.3995264498, 
    3059.84926316331, 
    3101.29928888572, 
    3121.75818816685, 
    3118.87626189301, 
    3196.72984270667, 
    3196.58785214621, 
    3140.11426193488, 
    3194.27228470368, 
    3242.2721838923, 
    3262.96465789327, 
    3297.80566248291, 
    3348.70705160651, 
    3378.60664970903, 
    3385.31401798131, 
    3383.19627292613, 
    3302.91301087063, 
    3326.46630085533, 
    3425.70909879532, 
    3589.35973357407, 
    3622.2018159527, 
    3543.67165433051, 
    3442.91012495132, 
    3372.88465217949, 
    3353.89210726396, 
    3442.20101396012, 
    3426.15148391248, 
    3406.15065085326, 
    3420.71660552436, 
    3587.83271368051, 
    3640.11971596856, 
    3643.51239125094, 
    3541.11643559626, 
    3349.67856206192, 
    3488.52520266396, 
    3539.99549668445, 
    3474.68042013551, 
    3425.03382271439, 
    3362.54893048401, 
    3435.97672726944, 
    3494.14398205922, 
    3356.92215828808, 
    3315.52831273752, 
    3198.90065253286, 
    3152.8273339568, 
    3115.40504829337, 
    3047.66250308298, 
    3000.34065300074, 
    3021.83743602508, 
    3092.2258326126, 
    3068.07259554813, 
    3025.85725460525, 
    2990.10010310319, 
    2970.775722929, 
    2898.11192093922, 
    2840.55786358389, 
    2805.2454707171, 
    2857.80483876077, 
    2763.23780490621, 
    2752.93767810663, 
    2759.62614546572, 
    2687.84723975149, 
    2608.51695643287, 
    2564.47696108435, 
    2400.36537371229, 
    2289.90146128691, 
    2311.00841999972, 
    2310.2756339256, 
    2135.12773754912, 
    1874.0681177874, 
    1732.56913178143, 
    1588.90197122725, 
    1422.32823592861, 
    1254.76882978469, 
    1087.69057113716, 
    959.089052032999, 
    923.328449496286, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    998.802722068279, 
    701.644338535775, 
    946.114299641018, 
    1168.87531025726, 
    2199.9780478282, 
    1916.9959294666, 
    1875.66205688186, 
    1841.89965105058, 
    1885.96939309532, 
    2175.01873198519, 
    2657.17375846181, 
    2969.87609284029, 
    2883.49061512766, 
    2705.66813099896, 
    2830.89116789233, 
    2855.33549999211, 
    3084.58236205981, 
    3119.53002638308, 
    3049.37744887685, 
    3063.6363787978, 
    3156.14167888613, 
    3101.97312069353, 
    3134.67063278169, 
    3246.89195884996, 
    3311.45834430519, 
    3328.85798974593, 
    3372.93959662643, 
    3399.32981653343, 
    3396.8443002114, 
    3401.00777781768, 
    3345.48364595625, 
    3323.84860460504, 
    3392.61143606953, 
    3533.83301195359, 
    3621.73323921658, 
    3576.76369452679, 
    3615.92303761329, 
    3384.0111389149, 
    3354.12314468025, 
    3384.18206457129, 
    3396.33952700205, 
    3487.29368317962, 
    3452.94453189716, 
    3463.68823900239, 
    3552.28878273744, 
    3615.53665912825, 
    3639.74483966033, 
    3577.85110843159, 
    3431.32688136272, 
    3446.97558369883, 
    3508.87324137319, 
    3462.70604048308, 
    3515.49831549262, 
    3361.57264861501, 
    3425.42662779559, 
    3464.42802505583, 
    3281.48997031941, 
    3171.5705193221, 
    3113.62105231238, 
    3061.04232995451, 
    3037.36352662695, 
    2962.01009975884, 
    2949.06415465557, 
    3003.48843688561, 
    3003.09529140694, 
    2993.05380399879, 
    2976.93004372106, 
    2942.86224845842, 
    2874.21182093368, 
    2792.64327919179, 
    2774.40407255294, 
    2779.98967902119, 
    2757.56330914563, 
    2640.46978121875, 
    2638.98942020243, 
    2632.22653758395, 
    2626.56511526319, 
    2592.37316248933, 
    2575.19390181792, 
    2368.4478329571, 
    2228.99844084175, 
    2126.49322508909, 
    2033.21478672942, 
    2128.21937233774, 
    1944.05214866042, 
    1735.25128572781, 
    1444.16081444052, 
    1371.31488801259, 
    1294.31771311618, 
    1119.86714868805, 
    524.480100844889, 
    761.96686802302, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1015.47691857508, 
    1565.75849384035, 
    1255.01181323545, 
    1260.53800655811, 
    1812.96388068967, 
    1099.83362851857, 
    1360.80946938186, 
    1604.10110269116, 
    1596.99270927005, 
    1733.12293289151, 
    2210.78680943101, 
    2523.81953626211, 
    2629.1279378322, 
    2820.24387078422, 
    2862.26510076539, 
    3016.51166465153, 
    3100.76971447612, 
    3018.20535820221, 
    3012.22572361767, 
    3051.3952844958, 
    3094.19762811275, 
    3085.86639503614, 
    3150.89895796043, 
    3288.50566253733, 
    3369.74258948653, 
    3346.50146922022, 
    3366.85484743476, 
    3412.3823418232, 
    3427.09305859389, 
    3356.55455619921, 
    3375.30854464384, 
    3367.72091749741, 
    3376.94470665793, 
    3454.25920533085, 
    3453.5125359901, 
    3496.82408652417, 
    3582.11626844155, 
    3398.38565699553, 
    3416.28591755517, 
    3399.29446801723, 
    3365.45252588024, 
    3545.0624753465, 
    3501.66546063425, 
    3465.00993549558, 
    3564.4251871419, 
    3397.61419424672, 
    3350.98941422805, 
    3464.7328591266, 
    3596.75649341761, 
    3527.74633206382, 
    3502.2944575625, 
    3334.26122472845, 
    3414.48468350116, 
    3373.44244357677, 
    3505.68579617258, 
    3427.23000646049, 
    3291.05278114895, 
    3067.23723196765, 
    3044.77872150185, 
    3016.40476861948, 
    2980.87564025974, 
    2889.21970282639, 
    2869.97196703052, 
    2898.75532279576, 
    2889.38063768554, 
    2908.4467629314, 
    2929.67538087176, 
    2917.03999999801, 
    2884.77423665023, 
    2829.68673057379, 
    2738.98163338081, 
    2715.11940554163, 
    2673.70224988176, 
    2587.29689678998, 
    2580.02353331236, 
    2580.40535570907, 
    2594.58416031601, 
    2567.93849208578, 
    2467.27678319807, 
    2397.53468283584, 
    2320.23678017029, 
    2233.65527310963, 
    2196.43769256374, 
    2220.64308737761, 
    1940.51262623624, 
    1578.42024885316, 
    1576.43535551905, 
    1415.01556711891, 
    1107.01128535798, 
    677.325051013744, 
    657.609301300825, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    767.822696264813, 
    1266.55662624847, 
    1505.21729125879, 
    1869.05436714982, 
    1158.44978333472, 
    884.62397065174, 
    863.978285977649, 
    1349.44984555908, 
    1319.33887097097, 
    1250.11720135672, 
    1712.18460205939, 
    2226.47246342779, 
    2817.87107873373, 
    2788.22261386755, 
    2749.62762755268, 
    2837.00198116208, 
    2977.0509629501, 
    2984.16156805927, 
    3019.21917419612, 
    3009.99176871732, 
    2949.74560587339, 
    3005.37577026268, 
    3118.71592936064, 
    3312.09818745351, 
    3447.84416715258, 
    3306.59463877055, 
    3256.87937443269, 
    3435.92741700213, 
    3423.83208114573, 
    3419.39934769451, 
    3333.97162476477, 
    3376.5560728573, 
    3376.70816355497, 
    3364.85182006515, 
    3556.22280868665, 
    3356.1408882129, 
    3408.27456857339, 
    3231.6229855456, 
    3258.58644818637, 
    3334.12423657811, 
    3333.52882360519, 
    3420.23465357652, 
    3494.52523598143, 
    3509.83838187765, 
    3437.88312590713, 
    3376.29825824655, 
    3336.33529841987, 
    3496.61850180237, 
    3575.9366002333, 
    3548.71099774311, 
    3420.13077150824, 
    3429.18215353096, 
    3424.66028867775, 
    3444.20374404337, 
    3501.09890120145, 
    3387.98554462371, 
    3294.45389347659, 
    3074.19959917879, 
    3045.11242254591, 
    3037.98068701636, 
    2909.19618518417, 
    2877.92452238754, 
    2831.12626994258, 
    2885.1411509587, 
    2813.42771452061, 
    2807.68553183001, 
    2888.60792385608, 
    2900.55637045934, 
    2857.79451636678, 
    2775.49067003843, 
    2827.80559531482, 
    2731.1445363764, 
    2579.05053575111, 
    2535.49115280592, 
    2549.73497101934, 
    2558.63025195697, 
    2495.29185658902, 
    2459.34976279054, 
    2446.81619333106, 
    2291.69819211042, 
    2271.66120355052, 
    2294.96002742536, 
    2198.56804051092, 
    2183.02571605828, 
    1981.17963607909, 
    1520.81833346249, 
    1519.43579979086, 
    1098.42531446434, 
    950.599519144118, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1074.9623660437, 
    827.806372449429, 
    645.841646693, 
    800.420137273776, 
    0, 
    0, 
    0, 
    1324.22076894677, 
    1640.16502430482, 
    1261.34283092024, 
    1545.24397019282, 
    1884.51457555217, 
    2194.15994189391, 
    2397.55839239656, 
    2565.65133533908, 
    2712.53140767814, 
    2971.35614638684, 
    3054.31436123808, 
    3088.41301993728, 
    3021.05630434978, 
    2915.29666173613, 
    2968.66560902832, 
    3192.33673574107, 
    3308.13470946113, 
    3454.80683408533, 
    3330.77101790922, 
    3256.27161367184, 
    3264.79379399418, 
    3374.49994046092, 
    3404.22234702788, 
    3289.99158337615, 
    3285.58731817762, 
    3350.30597208744, 
    3406.30139315061, 
    3498.99701881347, 
    3344.29765306245, 
    3052.5881251306, 
    3052.0416238191, 
    3067.76164013463, 
    3177.86741026987, 
    3287.79079408017, 
    3341.70393704821, 
    3377.1586767593, 
    3299.85259135502, 
    3200.90125620251, 
    3507.31631887489, 
    3335.56222148509, 
    3580.91311308994, 
    3474.65440360114, 
    3512.29588639611, 
    3363.37461937738, 
    3418.48864770048, 
    3412.33637907652, 
    3267.25018453857, 
    3351.6796846442, 
    3346.58374392645, 
    3236.17129568122, 
    3040.10762054547, 
    3016.75363578482, 
    2901.2282588579, 
    2785.20051988784, 
    2812.8197247128, 
    2773.15222506938, 
    2743.84783659492, 
    2772.06431234494, 
    2668.6138049725, 
    2729.86338949206, 
    2885.56943358012, 
    2867.13774526209, 
    2760.12848413203, 
    2680.09964949478, 
    2587.65060052684, 
    2498.66496971994, 
    2472.6813684787, 
    2474.94279536702, 
    2464.00076489608, 
    2423.76292113987, 
    2390.1209820818, 
    2353.32058307468, 
    2230.12902434782, 
    2205.30731572711, 
    2185.47388762865, 
    2110.40125469505, 
    2065.60137151481, 
    1981.81751208594, 
    1703.87584528512, 
    1393.88291829181, 
    998.533887674994, 
    1034.04898333161, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    944.670543879502, 
    860.156487877056, 
    0, 
    0, 
    0, 
    0, 
    0, 
    497.902117700483, 
    1185.66422485264, 
    1255.17410023979, 
    1541.54424570484, 
    1863.06585614588, 
    1970.90144054726, 
    2093.85579316286, 
    2424.46204760889, 
    2384.00330357164, 
    2769.74325619632, 
    3208.99129268543, 
    3269.70140288611, 
    2942.88312367663, 
    2739.22687355007, 
    2787.55911315015, 
    2955.52553271192, 
    3175.8176409897, 
    3297.9135276478, 
    3302.21099651246, 
    3293.09227234825, 
    3296.95322176454, 
    3397.50708361974, 
    3397.00676327081, 
    3397.03748176248, 
    3363.45487012257, 
    3286.49538276692, 
    3343.77963145427, 
    3384.14323314232, 
    3137.21600976822, 
    3308.21844620987, 
    3045.32347332443, 
    2893.37505145983, 
    2992.58011631595, 
    3119.13383274689, 
    3140.08682190198, 
    3030.73913520839, 
    2872.67960387896, 
    3064.17241759885, 
    3025.52828701323, 
    3156.51298479114, 
    3151.59093596568, 
    3235.87139099293, 
    3261.10705123685, 
    3175.57947124919, 
    3307.46403531614, 
    3167.23890412504, 
    2959.38142465403, 
    3087.69497489979, 
    3128.92228144936, 
    3043.33279717738, 
    2916.88913166093, 
    2919.52168111852, 
    2946.74013503917, 
    2787.33701129289, 
    2738.08361493618, 
    2730.170087893, 
    2660.04392690344, 
    2647.89903280047, 
    2633.53440784181, 
    2773.02755102257, 
    2837.48164576455, 
    2885.2837727874, 
    2719.95219354768, 
    2607.40583878644, 
    2503.65330895905, 
    2433.90957594704, 
    2430.44537581923, 
    2406.39616111003, 
    2362.73725364216, 
    2329.4629140254, 
    2317.14198906977, 
    2250.23633136804, 
    2147.45569120605, 
    2106.37814137764, 
    2023.41386403412, 
    1960.06573866903, 
    1859.61706727203, 
    1731.61735040848, 
    1850.80414528145, 
    1703.15346690792, 
    1522.66543217227, 
    1308.11943139789, 
    954.694898751642, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    984.684590409615, 
    1168.26539194608, 
    1533.65054777324, 
    1982.9739711832, 
    1354.88102394163, 
    1680.19369094981, 
    2260.99034693854, 
    2155.4486733418, 
    2846.82153970453, 
    3206.49943788774, 
    2979.55801116278, 
    2611.36349975258, 
    2401.91598952548, 
    2550.37474760415, 
    2686.16892012755, 
    2938.65570893609, 
    3214.47656622605, 
    3249.34286431011, 
    3335.19578391582, 
    3230.84090495375, 
    3357.90785818328, 
    3420.77231838082, 
    3387.07853183765, 
    3304.88979978442, 
    3288.77007395722, 
    3309.79123568042, 
    3441.46928226706, 
    3313.28539438549, 
    3169.50407958701, 
    3137.98443488729, 
    2906.73734784797, 
    2860.09893135469, 
    2779.6111133814, 
    2735.44655249024, 
    2781.47080789053, 
    2977.75978762722, 
    3230.77313634984, 
    2991.6655296922, 
    2778.98041313329, 
    2744.27373773734, 
    2814.45525951275, 
    3210.91268657694, 
    3144.2113541993, 
    3081.51121970621, 
    2870.29762167473, 
    2852.30038798731, 
    2891.32068733078, 
    3014.31790012563, 
    2946.41975581664, 
    2945.87032798569, 
    2986.61684303216, 
    3012.70743458484, 
    2912.33283037829, 
    2835.00634897175, 
    2785.96477931996, 
    2646.13063964543, 
    2590.54893239564, 
    2490.50300950997, 
    2563.96343675776, 
    2649.76815004526, 
    2733.85191313123, 
    2835.96951636935, 
    2622.23245879312, 
    2465.03890220927, 
    2415.59056154261, 
    2388.97018096684, 
    2330.81588832158, 
    2270.12954596532, 
    2126.90848676713, 
    2157.34511086008, 
    2124.32524675142, 
    2041.19594071006, 
    1949.69065089775, 
    1891.31433653735, 
    1794.95464836671, 
    1638.02114115503, 
    1558.7689537235, 
    1580.13432116937, 
    1740.22024484193, 
    1337.3156228671, 
    800.522997081661, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    788.120900618625, 
    1049.24041706163, 
    1350.16319386337, 
    1473.96452477921, 
    1610.34048043519, 
    1332.18073953392, 
    1293.07377117358, 
    1841.82149358423, 
    2159.78316081279, 
    2171.51728916798, 
    2491.58612460443, 
    2293.83563420723, 
    2237.31930339666, 
    2567.32483735073, 
    2727.01365587684, 
    2558.41069951807, 
    2768.62905633527, 
    2922.55121936327, 
    3176.01040194969, 
    3246.54044152528, 
    3198.34152424502, 
    3266.24787078619, 
    3265.36973694866, 
    3202.71247905981, 
    3212.78927845792, 
    3233.52054355778, 
    3245.03968492646, 
    3294.85911161997, 
    3285.01348120029, 
    3161.93726879887, 
    3013.00228375281, 
    2929.24927940131, 
    2967.25295467369, 
    2734.94702097839, 
    2440.23395168991, 
    2630.69389340305, 
    2828.79526736132, 
    2859.00346899562, 
    2875.59776128252, 
    2956.81093399931, 
    3106.69191784215, 
    3429.60580611576, 
    3345.10674229179, 
    3291.16538018823, 
    3007.1270771373, 
    2882.42339886815, 
    2772.21771744473, 
    2780.18064933069, 
    2772.24932438461, 
    2745.84270555384, 
    2743.75485575309, 
    2942.07598059577, 
    2999.34592727937, 
    2861.1212429218, 
    2906.88934056247, 
    2686.60331772904, 
    2647.59269258816, 
    2544.05664835958, 
    2354.84874153503, 
    2382.2781226011, 
    2423.58786461764, 
    2559.65763538256, 
    2673.22587536976, 
    2532.23132315865, 
    2440.64298325356, 
    2409.99316903555, 
    2355.15242196139, 
    2186.69617004277, 
    2105.27375242316, 
    2017.20282137471, 
    2007.73840846816, 
    1970.31710266471, 
    1893.69162062572, 
    1828.77589457596, 
    1746.60825420546, 
    1654.74312943238, 
    1489.48284513501, 
    1320.11970651572, 
    1278.45528849929, 
    1480.78783984349, 
    857.341952991517, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1174.11723438799, 
    574.518402166606, 
    994.27595631292, 
    1077.10070656687, 
    1640.01299720138, 
    1641.81917758631, 
    1198.48186799676, 
    1517.47740589733, 
    1675.84175100921, 
    2048.6452679149, 
    2421.18295490794, 
    1903.392187992, 
    1813.81648805787, 
    2598.17149638862, 
    2554.62947595653, 
    2177.90545661548, 
    2105.54436182804, 
    2590.55229676209, 
    2997.93645738017, 
    3111.67668160567, 
    3116.66951469906, 
    3218.29018378738, 
    3165.14488396223, 
    3165.43021764729, 
    3287.10468654058, 
    3099.30643610489, 
    3077.85892495797, 
    3214.40816957865, 
    3295.03859315054, 
    3215.5908511893, 
    3083.62079725256, 
    3004.93075626232, 
    3050.49565354863, 
    3013.34501743897, 
    2518.30751529159, 
    2795.98748955589, 
    2908.51692359197, 
    2657.13796401693, 
    2730.51150560663, 
    3012.90824715379, 
    3193.1314520831, 
    2830.58387062948, 
    2865.45966350557, 
    2853.69609616674, 
    2856.69002821238, 
    2925.41548321358, 
    2833.84204607554, 
    2686.53261027792, 
    2540.77104393348, 
    2589.85738430972, 
    2723.86262972863, 
    2887.1735576605, 
    2859.72361279658, 
    2569.99901302913, 
    2717.23996868929, 
    2864.87826802731, 
    2680.65721855258, 
    2704.97738660782, 
    2424.44793767562, 
    2296.81065903246, 
    2295.15405922482, 
    2247.09881775832, 
    2266.760773665, 
    2289.57798564089, 
    2334.24066508672, 
    2242.4001664128, 
    2163.34940024603, 
    2009.12650668803, 
    1987.13899061673, 
    1944.27639783561, 
    1933.92469562322, 
    1891.0964048347, 
    1768.14166595471, 
    1693.56862427799, 
    1608.41480026581, 
    1532.79143171384, 
    1387.31741127074, 
    1111.01431181547, 
    1127.37982292643, 
    876.078467028988, 
    1371.78811622039, 
    69.3978954424642, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    765.757680357693, 
    734.020923265824, 
    828.074465477041, 
    1126.49973298658, 
    1528.54883597838, 
    980.543419476799, 
    1071.02965430225, 
    1227.71375868396, 
    1619.50132865009, 
    1631.86635682685, 
    1879.38489136303, 
    1982.40362296175, 
    2572.18454474256, 
    2124.60511828554, 
    2155.91930201115, 
    2352.2642083821, 
    2626.78986513916, 
    2920.58664769285, 
    2980.67687244194, 
    3016.03989841437, 
    3054.9318582055, 
    3134.91674488616, 
    3086.23455238819, 
    3089.64846132958, 
    3062.94726197445, 
    2935.34335902104, 
    3055.5878636423, 
    3144.40591922133, 
    3202.32118298518, 
    3090.96937020774, 
    2762.729070141, 
    2963.18811280222, 
    2893.3504601841, 
    2707.76479564521, 
    2684.99948681452, 
    2489.32455419148, 
    2335.4986616488, 
    2335.60556566013, 
    2710.48771664626, 
    2883.60311669511, 
    2354.25217879587, 
    2425.21082139592, 
    2558.85521692554, 
    2592.082291814, 
    2929.8110199023, 
    2892.83543625961, 
    2628.92054325572, 
    2600.73896671599, 
    2710.91474833843, 
    2786.90927809208, 
    2846.1515732833, 
    2747.29250921261, 
    2658.75120180307, 
    2614.94572612458, 
    2701.87661843534, 
    2735.39855673314, 
    2397.34092641342, 
    2595.34037424715, 
    2273.27563864846, 
    2179.06736394557, 
    2155.92216007689, 
    2145.34499041737, 
    2107.98246278986, 
    2207.98420938515, 
    2338.96985967824, 
    2081.69159400404, 
    2044.80783628157, 
    1974.62269589149, 
    1947.97069096189, 
    1909.55090880303, 
    1823.13280865341, 
    1653.51479241139, 
    1537.06628871362, 
    1434.85612205055, 
    1188.76591298179, 
    1181.44317249062, 
    908.9967456127, 
    887.769673876361, 
    0, 
    0, 
    0, 
    3.82501220703125, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    830.42739181241, 
    815.397368016162, 
    956.425366172859, 
    865.194644233915, 
    1002.27231361998, 
    1043.41111255457, 
    1139.76392774609, 
    1205.80547146628, 
    1310.83935930463, 
    2091.56672462938, 
    2126.07849394993, 
    2129.8339636094, 
    1917.61041177616, 
    2176.0277945275, 
    2389.468625917, 
    2740.71306099343, 
    2913.90678375651, 
    2886.57058570063, 
    2884.50261747266, 
    2884.63687699207, 
    2913.12049217128, 
    2942.65585589233, 
    2845.37367447885, 
    2849.58560353623, 
    2914.99925026882, 
    2973.81691613048, 
    3057.92223486859, 
    3119.50424526189, 
    3125.12841625663, 
    2980.06893193258, 
    2951.41731718774, 
    2739.87171982614, 
    2531.59136548683, 
    2376.13401100675, 
    2251.44261509493, 
    2193.0736808992, 
    2332.72491662723, 
    2314.25609772196, 
    2472.5693777005, 
    2263.03142404281, 
    2398.09274433767, 
    2626.41250661682, 
    2856.44871438541, 
    2899.18400095805, 
    2837.37929173026, 
    2604.64355224782, 
    2632.25991099591, 
    2614.67439481073, 
    2651.69550877972, 
    2663.09897933284, 
    2532.1442782431, 
    2629.16558074488, 
    2532.11733971662, 
    2665.48519988198, 
    2847.64593238588, 
    2739.0390123658, 
    2392.12799135958, 
    2247.37193869582, 
    2218.04978547504, 
    2146.77708871167, 
    2026.70488663304, 
    1990.59171198008, 
    1977.74267263358, 
    1924.04073262403, 
    2057.07882424573, 
    1975.15812650937, 
    1955.96903845891, 
    1887.63455237789, 
    1796.35705392587, 
    1784.84181953551, 
    1538.25397075712, 
    1382.26154974847, 
    1257.74301006841, 
    1092.25095200464, 
    905.905085644944, 
    799.429924245896, 
    564.077768036345, 
    0, 
    0, 
    4.18057250976562, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    845.757994968337, 
    1095.19898575357, 
    1040.5030454413, 
    815.650366058583, 
    739.012044412202, 
    1370.96448530035, 
    1286.44503909714, 
    1643.00296492325, 
    2261.08361760582, 
    2096.47414352607, 
    2276.17759325286, 
    2227.37352803597, 
    2296.49110073434, 
    2417.18639063377, 
    2702.4989135225, 
    2756.77916111437, 
    2748.86758302569, 
    2763.74277102526, 
    2669.30828297481, 
    2639.54132157212, 
    2885.04339934583, 
    2833.96851628719, 
    2767.46839833349, 
    2799.61956520077, 
    2836.60539753603, 
    2829.45885490543, 
    2963.43021117785, 
    3057.48272872362, 
    2996.82750048494, 
    2914.33223543405, 
    2724.31266883768, 
    2546.88267979772, 
    2411.40680114153, 
    2340.70258630453, 
    2183.01213059591, 
    2055.96265460008, 
    2334.73616294476, 
    2628.87770399532, 
    2635.20857290997, 
    2775.23611276911, 
    2577.15596568331, 
    2616.51995524231, 
    2721.19255207279, 
    2785.82255158423, 
    2685.93687479601, 
    2672.81211697666, 
    2728.68857065838, 
    2617.26892259918, 
    2548.17311175409, 
    2622.70644073684, 
    2412.68011910237, 
    2336.6611567086, 
    2478.99373210542, 
    2432.74431983239, 
    2571.16940179924, 
    2678.33582937778, 
    2246.51311016825, 
    2372.58527798395, 
    2164.17162594976, 
    2119.77681337804, 
    1976.05175801233, 
    1978.26599019249, 
    1830.6798299485, 
    1937.07848687323, 
    1804.30072267607, 
    1805.41834338653, 
    1873.78616331401, 
    1774.80101247799, 
    1792.51118049165, 
    1560.80261720385, 
    1348.19358023352, 
    1114.21652937541, 
    1016.07753109341, 
    1105.11209840676, 
    855.256416749653, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1057.5371185721, 
    1409.63700656013, 
    1236.30607289644, 
    1014.25892401659, 
    675.960924767898, 
    565.203794731052, 
    778.045644419973, 
    957.880133203677, 
    1629.43788793094, 
    2390.74271141487, 
    2224.70369867201, 
    1597.872279103, 
    1816.12256442203, 
    2178.53028911603, 
    2462.21213134561, 
    2547.64579803854, 
    2562.35203218779, 
    2489.91336609649, 
    2542.92666740246, 
    2447.18770739947, 
    2466.49130100603, 
    2654.912588295, 
    2692.49897319043, 
    2678.37235716334, 
    2664.73572026569, 
    2785.30274990728, 
    2600.79594257682, 
    2503.14058093832, 
    2391.79345891189, 
    2817.36669970118, 
    2868.85356525083, 
    2408.18517523032, 
    2449.95514971566, 
    2369.88974180724, 
    2431.55836653251, 
    1971.346171286, 
    1989.81291660734, 
    2024.95775810378, 
    2240.55749990461, 
    2433.82814061486, 
    2305.33871744317, 
    2095.39883611933, 
    2302.55536014461, 
    2393.73911122887, 
    2636.38356323523, 
    2649.94669035694, 
    2410.90000681698, 
    2446.98287652864, 
    2365.88437073251, 
    2356.98918014795, 
    2490.60823443944, 
    2391.28375905881, 
    2327.24247157238, 
    2236.95741359469, 
    2403.84676122751, 
    2222.17769168115, 
    2377.65660887503, 
    2254.13969412092, 
    2048.17500590676, 
    1915.64923979731, 
    1937.5200187938, 
    1827.57046309772, 
    1960.47035089376, 
    1836.91675954795, 
    1875.48348073198, 
    1875.52399620152, 
    1879.14678504321, 
    1831.4147152014, 
    1843.76883216096, 
    1803.77225418586, 
    1560.30920292852, 
    1284.14412415812, 
    1142.41803317532, 
    1026.28207097067, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    837.297725928511, 
    1191.26550927253, 
    1107.44454424038, 
    2239.06188406356, 
    1278.19082592373, 
    665.581354732842, 
    960.256573678624, 
    1446.89296221694, 
    1890.58594884644, 
    2130.80692851249, 
    2188.9730770317, 
    2141.10205839404, 
    2233.85735813332, 
    2190.35858533879, 
    2225.96869102097, 
    2310.19048258226, 
    2426.55035534229, 
    2505.57387768515, 
    2555.32722643264, 
    2576.97737765501, 
    2589.91950958521, 
    2667.32240296366, 
    2188.49565909913, 
    2058.89491361232, 
    2169.37077070195, 
    2659.61980432881, 
    2298.17938915617, 
    2119.00430509279, 
    1793.9176458333, 
    1736.38427995396, 
    1647.76566753381, 
    1455.56283943556, 
    1546.3426972233, 
    1742.0173101626, 
    1736.91330139387, 
    1756.90259036733, 
    2008.96906305922, 
    1932.86695671295, 
    2143.9620387917, 
    2534.62595590237, 
    2719.8522382147, 
    2408.59622652688, 
    2251.96867550277, 
    2152.988737152, 
    2240.0639005611, 
    2247.8089400594, 
    2313.03881235284, 
    2139.6468894242, 
    2055.50250136383, 
    2255.91741175868, 
    2096.69140817824, 
    1962.30274415032, 
    2218.1685422701, 
    1967.31870520745, 
    2045.00748016719, 
    1948.97647423769, 
    2104.66211495638, 
    2138.32455024939, 
    1897.61724948435, 
    1952.3911975419, 
    1592.52210599142, 
    1938.70410959045, 
    1955.8344069915, 
    1947.45814682763, 
    1779.87174870235, 
    1620.44141710493, 
    1454.96482600793, 
    1403.1651100512, 
    874.337997500045, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1306.32561528111, 
    862.112012279028, 
    1629.05945193003, 
    1933.61551618211, 
    1112.03482174955, 
    0, 
    0, 
    857.00734612184, 
    1072.15798189605, 
    1536.56736347246, 
    2176.28549973895, 
    1979.12189005459, 
    1936.92743083638, 
    1801.34741455239, 
    1800.95497164647, 
    1930.59995784946, 
    2092.26688035518, 
    2165.74581810753, 
    2076.02696307475, 
    2133.96548292214, 
    2337.66869705232, 
    2182.24734278533, 
    2038.89081230768, 
    1931.52555959114, 
    1973.29838772831, 
    1875.87702965937, 
    2000.15340005787, 
    1922.0875098116, 
    1984.26770756734, 
    1727.97567446076, 
    1792.56421371803, 
    1353.41188509749, 
    1079.56140154917, 
    1241.46306413203, 
    1608.21846437633, 
    1279.03667438371, 
    1493.09623632935, 
    1665.59381201245, 
    1720.32402210849, 
    2080.46500154494, 
    2159.66332769029, 
    2348.27019465076, 
    2256.22863336323, 
    2217.99374711163, 
    1905.28956418165, 
    2168.42270239022, 
    2119.60714863192, 
    2137.2326497132, 
    1867.90300873834, 
    1700.22154252637, 
    2336.20556584706, 
    1866.60016667931, 
    1838.07950708432, 
    2001.61538622653, 
    2108.45943141037, 
    1928.46227855573, 
    1945.72142722482, 
    1743.93058309138, 
    2118.55887291702, 
    2090.39678486471, 
    2150.78760919762, 
    2058.54465950407, 
    2048.75808685662, 
    1916.56840974725, 
    1818.99481507592, 
    1644.84655098127, 
    1447.53192783731, 
    1324.15194399069, 
    1057.9573479145, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    985.829112058663, 
    489.526635406658, 
    0, 
    0, 
    865.458984167864, 
    951.582789174824, 
    958.261848684217, 
    1352.76001586533, 
    1578.53688765654, 
    1613.61747339298, 
    2142.97091293582, 
    1572.95454577575, 
    1521.08495389809, 
    1587.97957673328, 
    1725.13745429539, 
    1908.72106959548, 
    1646.2087154489, 
    1555.97058895216, 
    1826.92693173841, 
    1975.26817420828, 
    1675.03435471406, 
    1191.00828218082, 
    1538.43375189882, 
    1486.26839649642, 
    1646.84697181188, 
    1651.17874864586, 
    1751.3886826456, 
    1939.81281545586, 
    1146.67062843527, 
    829.321434149461, 
    911.713599574694, 
    869.873409464896, 
    755.7456419258, 
    930.464291555814, 
    1336.38114742748, 
    1484.10723339833, 
    1463.18355536229, 
    1550.11238175006, 
    1706.31680814178, 
    2025.30562156317, 
    2150.98001120049, 
    2016.29767154787, 
    1789.46955233123, 
    1950.71152124722, 
    2076.856632497, 
    2043.71562413745, 
    1608.96125222255, 
    1584.34111513212, 
    1763.65853554933, 
    1382.92534485788, 
    1349.2510421581, 
    1755.11138903718, 
    1882.38558793655, 
    1637.55404456642, 
    1488.00969179264, 
    1706.12356297091, 
    1859.62911244698, 
    2051.99525474514, 
    2084.65403584158, 
    2057.65442416464, 
    2074.74993099083, 
    1974.71105057567, 
    1839.60386834919, 
    1609.02866745463, 
    1382.5277530883, 
    1067.69265219409, 
    285.081366215127, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1093.93055295776, 
    0, 
    0, 
    780.153602689339, 
    887.089152016976, 
    782.695736280625, 
    920.416603442198, 
    1076.48034119542, 
    1034.87604249228, 
    1260.60244491449, 
    1619.43317894805, 
    1660.10689349139, 
    1634.40545728192, 
    1292.43699745149, 
    1418.16160095166, 
    1979.28205729799, 
    1593.84909868986, 
    1132.59478158628, 
    1104.49512743047, 
    1932.10376805573, 
    1520.49069551839, 
    1404.9104142634, 
    1536.74944193916, 
    1402.45295436326, 
    1834.08153575543, 
    1292.06992608772, 
    1314.33653839354, 
    1127.67902497009, 
    876.965664710464, 
    0, 
    0, 
    0, 
    0, 
    312.01606855336, 
    943.827257885296, 
    1610.7150524511, 
    1442.09233325117, 
    1571.26907104114, 
    1867.18356470243, 
    2044.35022396634, 
    1996.90398143635, 
    1932.31125904992, 
    2073.38514343251, 
    1943.95856184116, 
    1919.71463086001, 
    1172.74807490974, 
    809.446721858487, 
    1045.12741820081, 
    1605.54211657043, 
    1151.35536167187, 
    970.997057475146, 
    1480.75732729025, 
    1777.2036613266, 
    1883.26070433056, 
    1759.42754301948, 
    1611.1746495531, 
    1362.15848743701, 
    1458.17776574159, 
    1653.6515309237, 
    1606.38407169366, 
    1699.54987663687, 
    1826.45990368164, 
    1759.84296967586, 
    1726.35604012752, 
    1474.53306990516, 
    1067.8288816166, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    741.594569075701, 
    2037.86767059278, 
    2072.76894036102, 
    1500.89815701933, 
    1083.3919195766, 
    1185.81124871796, 
    860.364415266486, 
    892.22168779019, 
    1135.00462661981, 
    1129.97074513647, 
    1373.86287280905, 
    1514.16162448139, 
    1047.07302537156, 
    932.590877320368, 
    1458.43583261018, 
    932.052539425107, 
    1066.64335766532, 
    1217.02959535621, 
    1416.7638950256, 
    1251.60729408375, 
    1276.29496060739, 
    1161.8721981382, 
    1237.75962789774, 
    1257.65535570366, 
    1238.56441951029, 
    520.398893195919, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    883.752356004429, 
    1061.62706131705, 
    1267.3216485385, 
    2136.3229459417, 
    1537.39036579232, 
    2083.65645196749, 
    2166.65389453323, 
    1953.74222482327, 
    1555.45423315636, 
    1377.79228622691, 
    1009.41302900425, 
    966.243675587782, 
    0, 
    474.783454774249, 
    552.054182115533, 
    933.481817652518, 
    618.535656031168, 
    730.804221040376, 
    993.369517934416, 
    1388.45909200336, 
    1404.8425165905, 
    957.182974684393, 
    1031.13811243756, 
    856.209166750717, 
    881.274528444706, 
    701.095910927694, 
    1143.96879343949, 
    1546.81006185485, 
    1775.91769493873, 
    1507.26224818051, 
    1597.20167359909, 
    1161.35696315088, 
    0, 
    0, 
    0, 
    0, 
    0, 
    906.574194190222, 
    544.803947489153, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    918.276312820674, 
    1812.89314583922, 
    1055.27789172318, 
    847.917023203251, 
    867.122529677526, 
    0, 
    0, 
    0, 
    733.314883432292, 
    587.106685983049, 
    840.797670831758, 
    1483.82080684213, 
    1181.66477073962, 
    1158.52200587704, 
    1355.35951371161, 
    1916.19707382072, 
    983.015094153485, 
    1122.60517088253, 
    1227.13902093786, 
    836.755328582044, 
    1269.99398568927, 
    1962.7102229394, 
    840.891046371454, 
    834.37550244309, 
    1171.0254622879, 
    1256.70588613553, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    878.137596281293, 
    993.739848074278, 
    1062.64245122095, 
    1307.9993490627, 
    1662.08249713511, 
    1857.52031389407, 
    1607.9386098089, 
    1725.63324162767, 
    2089.97243367305, 
    1258.08261591952, 
    618.702177289142, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    952.151237280224, 
    1591.38147861121, 
    1295.07269629813, 
    808.423827630654, 
    790.008444064386, 
    1088.28824818552, 
    1128.99500641512, 
    737.255438996352, 
    820.043406962416, 
    1634.71465495157, 
    1556.62163762755, 
    779.130902473013, 
    39.9435036783521, 
    527.569758526009, 
    41.8680305480957, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    726.892582959974, 
    602.267872689934, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    913.232462294822, 
    921.86053919245, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    1035.14018398124, 
    1314.55419583033, 
    1334.56619526627, 
    658.731909096726, 
    1015.74437353782, 
    983.467033827534, 
    703.454694124254, 
    0, 
    1251.84321965091, 
    955.862093885278, 
    1650.57966745494, 
    0, 
    701.985312884444, 
    922.767869226506, 
    814.957996607293, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    867.608478390918, 
    762.666730509882, 
    1236.84654361045, 
    1553.70600241615, 
    1315.63954338103, 
    1866.77226134251, 
    1701.99234961333, 
    1193.70963576074, 
    1057.55250584341, 
    859.078101272472, 
    0, 
    0, 
    0, 
    0, 
    0, 
    776.22329283757, 
    1369.96718448734, 
    1756.83718156623, 
    1099.1188340274, 
    810.195103179266, 
    0, 
    0, 
    0, 
    0, 
    800.388873705543, 
    1137.78695761873, 
    1330.41559720837, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    863.228355798299, 
    673.879051342675, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    823.159977452749, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    798.347549006236, 
    0, 
    0, 
    1467.59178688452, 
    1282.03662077585, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    662.580838581032, 
    1197.78686063647, 
    1260.59112583318, 
    1316.41643444217, 
    1477.39340978039, 
    1377.88566001779, 
    1481.54074308928, 
    1509.99204231875, 
    1736.92629580389, 
    1253.18651975699, 
    0, 
    0, 
    0, 
    0, 
    815.295330764737, 
    1484.61880782361, 
    1357.40834372074, 
    1257.05212354761, 
    1181.60823436977, 
    0, 
    0, 
    0, 
    0, 
    0, 
    680.602602694617, 
    714.786901197933, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    721.872001523953, 
    752.503697462655, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    601.834621555847, 
    1384.42397156109, 
    1565.51648336493, 
    1224.50133473474, 
    1177.46223390534, 
    1019.44707905895, 
    849.362368597881, 
    1318.4173531862, 
    1170.68299695016, 
    960.788011506674, 
    848.103718572769, 
    0, 
    20.0582370758057, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    60.9751014709473, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    929.041771643469, 
    1228.02552648466, 
    961.234406031434, 
    735.076650117795, 
    1013.63643202855, 
    515.756599710857, 
    538.510313180597, 
    921.31526192845, 
    272.68545835015, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    3.9305419921875, 
    0, 
    0, 
    10.3054335954783, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    18.1499633789062, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0,
  0, 0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 
    0, 0 ;

 topg =
  
    -3411.75952148438, 
    -3403.677734375, 
    -3461.13452148438, 
    -3417.931640625, 
    -3381.58227539062, 
    -3377.28491210938, 
    -3355.4736328125, 
    -3313.7216796875, 
    -3289.90551757812, 
    -3280.86303710938, 
    -3243.09936523438, 
    -3204.67895507812, 
    -3143.73657226562, 
    -3107.47338867188, 
    -3051.24829101562, 
    -2993.43408203125, 
    -2951.60424804688, 
    -2910.73559570312, 
    -2909.83422851562, 
    -2834.33325195312, 
    -2801.56982421875, 
    -2716.8232421875, 
    -2626.19116210938, 
    -2523.56958007812, 
    -2471.64013671875, 
    -2273.42993164062, 
    -1777.63012695312, 
    -1495.51086425781, 
    -1194.65209960938, 
    -1097.048828125, 
    -1130.42578125, 
    -1191.27319335938, 
    -1205.81115722656, 
    -1129.3974609375, 
    -1034.05749511719, 
    -940.295471191406, 
    -890.219421386719, 
    -879.535217285156, 
    -829.042663574219, 
    -779.467346191406, 
    -742.308776855469, 
    -708.685729980469, 
    -668.054931640625, 
    -625.153625488281, 
    -590.06005859375, 
    -592.140197753906, 
    -619.106201171875, 
    -652.474487304688, 
    -674.548583984375, 
    -729.968505859375, 
    -815.505981445312, 
    -739.854248046875, 
    -493.187713623047, 
    -244.056594848633, 
    -269.6826171875, 
    -314.234466552734, 
    -399.702850341797, 
    -326.203155517578, 
    -313.745330810547, 
    -316.535278320312, 
    -346.998168945312, 
    -488.744171142578, 
    -998.799621582031, 
    -1412.86291503906, 
    -1470.72412109375, 
    -1414.72216796875, 
    -1275.51318359375, 
    -919.049865722656, 
    -640.533447265625, 
    -625.350341796875, 
    -812.410827636719, 
    -921.275573730469, 
    -1041.62561035156, 
    -1377.69445800781, 
    -1705.408203125, 
    -1869.96813964844, 
    -1997.81567382812, 
    -2094.6796875, 
    -2159.44506835938, 
    -2191.06176757812, 
    -2194.96264648438, 
    -2224.9111328125, 
    -2215.33447265625, 
    -2201.00390625, 
    -2181.07250976562, 
    -2179.62890625, 
    -2248.85400390625, 
    -2149.73120117188, 
    -2184.01611328125, 
    -2226.986328125, 
    -2315.95239257812, 
    -2286.14672851562, 
    -2259.7451171875, 
    -2229.08935546875, 
    -2203.47045898438, 
    -2153.80932617188, 
    -2066.21557617188, 
    -1837.90270996094, 
    -1408.60498046875, 
    -790.149719238281, 
    -651.296752929688, 
    -577.519226074219, 
    -536.570068359375, 
    -525.099243164062, 
    -565.119995117188, 
    -587.210876464844, 
    -619.664916992188, 
    -651.612243652344, 
    -504.728302001953, 
    -267.361022949219, 
    -172.372375488281, 
    -200.293365478516, 
    -461.326019287109, 
    -598.764465332031, 
    -698.946960449219, 
    -669.763549804688, 
    -645.16064453125, 
    -531.925598144531, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -463.658996582031, 
    -200, 
    -207.519866943359, 
    -200, 
    -2300, 
    -2300, 
    -2300,
  
    -3413.40087890625, 
    -3438.47216796875, 
    -3472.67822265625, 
    -3395.91821289062, 
    -3372.9892578125, 
    -3371.98681640625, 
    -3334.78295898438, 
    -3311.78125, 
    -3291.96508789062, 
    -3271.64331054688, 
    -3254.44775390625, 
    -3244.61303710938, 
    -3163.4482421875, 
    -3120.32690429688, 
    -3057.60473632812, 
    -3016.1396484375, 
    -2979.93676757812, 
    -2925.00756835938, 
    -2898.43359375, 
    -2854.51416015625, 
    -2824.58959960938, 
    -2756.48413085938, 
    -2629.25512695312, 
    -2507.57348632812, 
    -2451.21118164062, 
    -1804.30712890625, 
    -1646.02136230469, 
    -1274.56848144531, 
    -1128.15832519531, 
    -1092.0400390625, 
    -1108.70373535156, 
    -1149.54663085938, 
    -1103.310546875, 
    -1019.68829345703, 
    -847.347412109375, 
    -504.027130126953, 
    -546.885131835938, 
    -759.495178222656, 
    -778.568298339844, 
    -766.281066894531, 
    -734.598205566406, 
    -676.947875976562, 
    -604.934387207031, 
    -432.078674316406, 
    -226.905212402344, 
    -204.51025390625, 
    -376.254852294922, 
    -490.843353271484, 
    -575.288146972656, 
    -644.702758789062, 
    -612.875549316406, 
    -402.4140625, 
    -217.456436157227, 
    -212.981674194336, 
    -275.520477294922, 
    -322.629974365234, 
    -351.164886474609, 
    -340.835052490234, 
    -332.508819580078, 
    -344.996459960938, 
    -328.606628417969, 
    -337.092102050781, 
    -518.286315917969, 
    -935.928344726562, 
    -1253.80603027344, 
    -1164.74108886719, 
    -838.137084960938, 
    -427.837677001953, 
    -488.596038818359, 
    -524.984802246094, 
    -677.563171386719, 
    -709.115905761719, 
    -833.987487792969, 
    -1029.45190429688, 
    -1312.69580078125, 
    -1632.35302734375, 
    -1773.18566894531, 
    -1920.4912109375, 
    -2008.10791015625, 
    -2108.21533203125, 
    -2112.30688476562, 
    -2121.99584960938, 
    -2125.69555664062, 
    -2119.98486328125, 
    -2095.25561523438, 
    -2037.86364746094, 
    -2033.67895507812, 
    -1913.40588378906, 
    -1854.705078125, 
    -1948.60620117188, 
    -2054.60913085938, 
    -2070.00244140625, 
    -2070.51098632812, 
    -2225.78784179688, 
    -2212.28491210938, 
    -2207.6376953125, 
    -1994.08581542969, 
    -1458.87084960938, 
    -699.539245605469, 
    -470.33447265625, 
    -421.278686523438, 
    -462.302703857422, 
    -486.099517822266, 
    -457.916687011719, 
    -448.721557617188, 
    -487.284118652344, 
    -298.429168701172, 
    -230.528106689453, 
    -449.495880126953, 
    -717.349304199219, 
    -831.015258789062, 
    -506.321990966797, 
    -308.888275146484, 
    -333.002258300781, 
    -306.084747314453, 
    -381.34521484375, 
    -670.432189941406, 
    -640.883361816406, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -202.870727539062, 
    -646.013061523438, 
    -677.536010742188, 
    -747.549011230469, 
    -734.746520996094, 
    -2300, 
    -2300,
  
    -3460.6875, 
    -3436.32983398438, 
    -3411.95434570312, 
    -3390.12255859375, 
    -3391.33959960938, 
    -3371.19458007812, 
    -3325.27294921875, 
    -3305.92797851562, 
    -3281.88110351562, 
    -3259.37426757812, 
    -3262.18969726562, 
    -3198.80053710938, 
    -3142.82568359375, 
    -3096.45068359375, 
    -3095.98828125, 
    -3051.48706054688, 
    -3002.541015625, 
    -2936.67407226562, 
    -2893.9091796875, 
    -2865.86401367188, 
    -2844.20971679688, 
    -2745.78759765625, 
    -2624.60766601562, 
    -2491.86010742188, 
    -2397.13916015625, 
    -1686.47875976562, 
    -1394.2802734375, 
    -1153.81958007812, 
    -1038.96862792969, 
    -1059.80212402344, 
    -1215.0263671875, 
    -1078.70581054688, 
    -984.425903320312, 
    -726.271606445312, 
    -268.134155273438, 
    -271.50244140625, 
    -293.224182128906, 
    -503.169036865234, 
    -640.347778320312, 
    -590.735168457031, 
    -533.891906738281, 
    -382.680053710938, 
    -220.713027954102, 
    -157.792572021484, 
    -203.958602905273, 
    -169.991592407227, 
    -170.429870605469, 
    -167.497604370117, 
    -212.767349243164, 
    -266.735778808594, 
    -271.28125, 
    -206.123474121094, 
    -200.364776611328, 
    -210.975311279297, 
    -235.542251586914, 
    -297.180358886719, 
    -385.621490478516, 
    -329.973571777344, 
    -343.571655273438, 
    -301.097961425781, 
    -300.500213623047, 
    -307.367034912109, 
    -311.4580078125, 
    -426.729309082031, 
    -500.503356933594, 
    -567.268249511719, 
    -405.028350830078, 
    -342.394226074219, 
    -411.328399658203, 
    -514.920776367188, 
    -639.136108398438, 
    -614.61083984375, 
    -627.077270507812, 
    -782.881652832031, 
    -962.224792480469, 
    -1171.69982910156, 
    -1473.95202636719, 
    -1642.15478515625, 
    -1800.16540527344, 
    -1886.16687011719, 
    -1931.09069824219, 
    -1788.30786132812, 
    -1811.73840332031, 
    -1915.11328125, 
    -1978.65600585938, 
    -1867.86157226562, 
    -1578.74670410156, 
    -828.231140136719, 
    -672.350524902344, 
    -735.939453125, 
    -1108.88305664062, 
    -1387.67272949219, 
    -1611.97424316406, 
    -1953.73583984375, 
    -1929.53356933594, 
    -1618.36779785156, 
    -1383.39489746094, 
    -778.169616699219, 
    -506.643188476562, 
    -428.841857910156, 
    -387.821014404297, 
    -379.539703369141, 
    -317.797943115234, 
    -315.617370605469, 
    -154.959014892578, 
    -117.034729003906, 
    -83.5130767822266, 
    -54.386100769043, 
    -170.152694702148, 
    -124.344093322754, 
    -228.452072143555, 
    -868.977478027344, 
    -248.554794311523, 
    -74.8536148071289, 
    -172.778472900391, 
    -260.138427734375, 
    -562.851745605469, 
    -675.407958984375, 
    -507.712585449219, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200.677642822266, 
    -200, 
    -200, 
    -200, 
    -215.683441162109, 
    -524.49072265625, 
    -483.828216552734, 
    -266.461395263672, 
    -200, 
    -200, 
    -804.895263671875, 
    -2300,
  
    -3477.32177734375, 
    -3421.81127929688, 
    -3412.78344726562, 
    -3401.52978515625, 
    -3382.23974609375, 
    -3359.86303710938, 
    -3329.18237304688, 
    -3308.12939453125, 
    -3278.40161132812, 
    -3245.99658203125, 
    -3207.3427734375, 
    -3129.1103515625, 
    -3076.63818359375, 
    -3042.29516601562, 
    -3009.375, 
    -2990.36059570312, 
    -2997.87475585938, 
    -2937.40014648438, 
    -2868.60693359375, 
    -2833.56176757812, 
    -2806.03979492188, 
    -2760.90502929688, 
    -2621.36743164062, 
    -2434.49633789062, 
    -2282.18310546875, 
    -1590.4140625, 
    -1345.93115234375, 
    -1236.22863769531, 
    -1160.28735351562, 
    -1308.35852050781, 
    -1291.19458007812, 
    -1073.21630859375, 
    -734.719482421875, 
    -235.820373535156, 
    -160.536254882812, 
    -162.541030883789, 
    -201.101806640625, 
    -185.879684448242, 
    -151.720520019531, 
    -123.931045532227, 
    -108.605323791504, 
    -132.880294799805, 
    -116.158210754395, 
    -130.867431640625, 
    -202.788131713867, 
    -198.319351196289, 
    -178.987762451172, 
    -147.742599487305, 
    -135.411346435547, 
    -113.957305908203, 
    -121.897354125977, 
    -132.027969360352, 
    -146.666046142578, 
    -181.876190185547, 
    -179.845962524414, 
    -215.224487304688, 
    -321.175872802734, 
    -357.646270751953, 
    -348.449249267578, 
    -322.298828125, 
    -299.441986083984, 
    -297.530975341797, 
    -299.502563476562, 
    -287.080810546875, 
    -307.480072021484, 
    -319.824188232422, 
    -293.251129150391, 
    -293.051239013672, 
    -327.714477539062, 
    -460.385528564453, 
    -599.86865234375, 
    -524.479125976562, 
    -403.691650390625, 
    -458.932861328125, 
    -636.453125, 
    -801.728942871094, 
    -1000.43701171875, 
    -1197.4169921875, 
    -1414.62548828125, 
    -1513.15026855469, 
    -1367.58422851562, 
    -1030.79626464844, 
    -1027.23413085938, 
    -1341.84973144531, 
    -1668.20153808594, 
    -1511.69702148438, 
    -803.161376953125, 
    -482.382385253906, 
    -591.652282714844, 
    -700.183837890625, 
    -782.228271484375, 
    -808.056518554688, 
    -938.963012695312, 
    -1298.43249511719, 
    -1224.92224121094, 
    -690.956481933594, 
    -513.611145019531, 
    -380.283477783203, 
    -318.711273193359, 
    -354.885131835938, 
    -383.720031738281, 
    -412.365936279297, 
    -196.685836791992, 
    -119.97297668457, 
    369.036102294922, 
    327.938903808594, 
    252.857925415039, 
    -33.7421951293945, 
    198.841262817383, 
    528.541687011719, 
    714.519470214844, 
    -712.6376953125, 
    86.1533966064453, 
    -106.387176513672, 
    -107.570686340332, 
    -118.771697998047, 
    -246.952011108398, 
    -652.446960449219, 
    -560.2822265625, 
    -298.085021972656, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -204.359344482422, 
    -238.269714355469, 
    -421.029418945312, 
    -705.031005859375, 
    -221.518768310547, 
    -200, 
    -200, 
    -200, 
    -201.572280883789, 
    -200, 
    -1483.33337402344,
  
    -3441.25366210938, 
    -3454.2802734375, 
    -3416.39990234375, 
    -3396.92846679688, 
    -3375.26342773438, 
    -3351.21826171875, 
    -3329.15502929688, 
    -3300.357421875, 
    -3282.26708984375, 
    -3215.60473632812, 
    -3170.15844726562, 
    -3103.11328125, 
    -3049.45776367188, 
    -3005.54931640625, 
    -2989.42895507812, 
    -2955.626953125, 
    -2950.39233398438, 
    -2912.07788085938, 
    -2864.80859375, 
    -2809.80615234375, 
    -2763.97924804688, 
    -2722.80786132812, 
    -2643.78369140625, 
    -2469.06469726562, 
    -2387.17944335938, 
    -2301.42944335938, 
    -2073.15551757812, 
    -1872.83203125, 
    -1528.29211425781, 
    -1266.95239257812, 
    -1048.54541015625, 
    -271.038787841797, 
    -286.158508300781, 
    -117.162590026855, 
    -132.933883666992, 
    -142.442749023438, 
    -121.231826782227, 
    -107.67456817627, 
    -109.048248291016, 
    -105.919486999512, 
    -109.18433380127, 
    -131.113708496094, 
    -105.368865966797, 
    -109.407836914062, 
    -151.931121826172, 
    -230.192031860352, 
    -141.573333740234, 
    -105.06388092041, 
    -91.1327819824219, 
    -110.801391601562, 
    -98.7336959838867, 
    -105.432731628418, 
    -129.580215454102, 
    -129.979354858398, 
    -148.28776550293, 
    -161.335586547852, 
    -315.576324462891, 
    -389.303192138672, 
    -340.132476806641, 
    -302.560638427734, 
    -275.387359619141, 
    -242.0146484375, 
    -284.465026855469, 
    -271.917907714844, 
    -268.067657470703, 
    -283.827209472656, 
    -328.593994140625, 
    -347.268218994141, 
    -330.123229980469, 
    -452.574035644531, 
    -589.276123046875, 
    -487.310516357422, 
    -376.640045166016, 
    -352.853149414062, 
    -420.773529052734, 
    -459.967559814453, 
    -576.660400390625, 
    -687.67724609375, 
    -943.192321777344, 
    -1024.05920410156, 
    -691.483032226562, 
    -690.270080566406, 
    -712.260925292969, 
    -833.119445800781, 
    -871.330017089844, 
    -440.048370361328, 
    -416.411895751953, 
    -474.858642578125, 
    -568.287963867188, 
    -672.050170898438, 
    -725.413024902344, 
    -756.540588378906, 
    -539.874694824219, 
    -652.971923828125, 
    -507.505279541016, 
    -365.607818603516, 
    -333.662811279297, 
    -313.765106201172, 
    -246.855743408203, 
    -199.628021240234, 
    -459.285766601562, 
    -551.136596679688, 
    -156.597274780273, 
    360.447235107422, 
    349.991668701172, 
    513.033325195312, 
    168.914947509766, 
    280.082000732422, 
    541.436096191406, 
    284.380554199219, 
    819.860168457031, 
    -644.933471679688, 
    63.2493629455566, 
    -66.2151184082031, 
    -109.501136779785, 
    109.598861694336, 
    131.817489624023, 
    -288.970306396484, 
    -486.975219726562, 
    -296.655609130859, 
    -200, 
    -200, 
    -213.249298095703, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -285.071960449219, 
    -327.683715820312, 
    -200, 
    -200, 
    -200, 
    -200.991256713867, 
    -200, 
    -200, 
    -200,
  
    -3454.30834960938, 
    -3433.26806640625, 
    -3413.54809570312, 
    -3398.87280273438, 
    -3391.30249023438, 
    -3387.8330078125, 
    -3312.53247070312, 
    -3272.53491210938, 
    -3208.16772460938, 
    -3189.484375, 
    -3130.9794921875, 
    -3081.3994140625, 
    -3004.62548828125, 
    -2981.783203125, 
    -2945.96997070312, 
    -2922.92407226562, 
    -2894.427734375, 
    -2879.0498046875, 
    -2814.19458007812, 
    -2752.18212890625, 
    -2724.57275390625, 
    -2671.50854492188, 
    -2565.58325195312, 
    -2446.05102539062, 
    -1994.96264648438, 
    -1589.27062988281, 
    -1390.08935546875, 
    -591.647338867188, 
    -373.767700195312, 
    -139.677627563477, 
    -88.1795883178711, 
    -200.867279052734, 
    -365.357360839844, 
    -119.696754455566, 
    -149.170013427734, 
    -142.704071044922, 
    -90.3420257568359, 
    -78.2760391235352, 
    -123.530227661133, 
    -105.66650390625, 
    -107.292434692383, 
    -97.848014831543, 
    -97.3846740722656, 
    -81.183723449707, 
    -64.7797698974609, 
    -340.008087158203, 
    -83.8657608032227, 
    -58.1435432434082, 
    -83.2720413208008, 
    -74.0015335083008, 
    -56.7941703796387, 
    -61.0527877807617, 
    -73.0999450683594, 
    -96.458137512207, 
    -107.471214294434, 
    -141.742904663086, 
    -431.769348144531, 
    -448.947479248047, 
    -343.85302734375, 
    -234.568588256836, 
    -200.554443359375, 
    -210.660430908203, 
    -189.679611206055, 
    -222.276336669922, 
    -217.500305175781, 
    -227.919174194336, 
    -283.079345703125, 
    -317.790679931641, 
    -360.0087890625, 
    -493.306549072266, 
    -506.104034423828, 
    -420.235900878906, 
    -393.428405761719, 
    -339.936920166016, 
    -333.261749267578, 
    -398.916534423828, 
    -439.613372802734, 
    -463.736389160156, 
    -444.494354248047, 
    -395.966827392578, 
    -468.703857421875, 
    -604.639587402344, 
    -690.307312011719, 
    -405.225891113281, 
    -457.037292480469, 
    -354.728240966797, 
    -406.424774169922, 
    -493.427764892578, 
    -573.046264648438, 
    -655.879821777344, 
    -665.891357421875, 
    -678.399658203125, 
    -289.592681884766, 
    -411.972961425781, 
    -302.435852050781, 
    -266.3984375, 
    -251.654922485352, 
    -213.869262695312, 
    -207.317825317383, 
    -379.558898925781, 
    -551.751586914062, 
    -688.29736328125, 
    -444.947601318359, 
    209.575653076172, 
    303.416656494141, 
    554.358337402344, 
    302.391662597656, 
    419.822235107422, 
    716.600036621094, 
    905.966674804688, 
    -287.778991699219, 
    -307.135284423828, 
    239.833190917969, 
    57.0292816162109, 
    430.024993896484, 
    712.388916015625, 
    854.488891601562, 
    322.127777099609, 
    -373.234832763672, 
    -392.351898193359, 
    -295.606048583984, 
    -367.178161621094, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -502.454986572266, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3450.09106445312, 
    -3417.1337890625, 
    -3394.46533203125, 
    -3397.98120117188, 
    -3387.09497070312, 
    -3352.85913085938, 
    -3270.45263671875, 
    -3202.45043945312, 
    -3150.66479492188, 
    -3092.27026367188, 
    -3067.7626953125, 
    -3006.17553710938, 
    -2981.10864257812, 
    -2968.4501953125, 
    -2923.72778320312, 
    -2908.96533203125, 
    -2844.09521484375, 
    -2773.9228515625, 
    -2723.4072265625, 
    -2633.9921875, 
    -2524.88623046875, 
    -2450.04345703125, 
    -2140.70556640625, 
    -1658.98083496094, 
    -552.474792480469, 
    -156.951644897461, 
    -93.5471496582031, 
    -104.515151977539, 
    -200.413421630859, 
    -39.7728462219238, 
    -45.0646705627441, 
    -64.9928512573242, 
    -220.210006713867, 
    -471.001892089844, 
    -433.426391601562, 
    -362.815734863281, 
    -154.065093994141, 
    -108.45027923584, 
    -138.494857788086, 
    -126.328216552734, 
    -165.803375244141, 
    -101.32625579834, 
    -76.4336395263672, 
    -53.5571708679199, 
    -49.9369201660156, 
    -147.27099609375, 
    -205.131576538086, 
    -37.8181266784668, 
    -64.9956817626953, 
    -50.8311996459961, 
    -49.9953880310059, 
    -49.9191246032715, 
    -42.724479675293, 
    -49.4221229553223, 
    -63.3225555419922, 
    -152.983337402344, 
    -505.612487792969, 
    -416.928649902344, 
    -264.460754394531, 
    -151.105804443359, 
    -148.331436157227, 
    -191.103912353516, 
    -194.320419311523, 
    -227.256011962891, 
    -198.628662109375, 
    -175.768981933594, 
    -239.236404418945, 
    -313.578826904297, 
    -390.147766113281, 
    -461.15576171875, 
    -491.590545654297, 
    -376.378540039062, 
    -324.349700927734, 
    -278.837707519531, 
    -303.253112792969, 
    -335.796539306641, 
    -370.174926757812, 
    -393.011840820312, 
    -305.327117919922, 
    -285.149780273438, 
    -350.005950927734, 
    -527.337768554688, 
    -686.015502929688, 
    -555.277709960938, 
    -354.934661865234, 
    -388.605224609375, 
    -383.454071044922, 
    -471.803771972656, 
    -544.57763671875, 
    -604.661560058594, 
    -613.464721679688, 
    -686.765258789062, 
    -401.497924804688, 
    -401.345001220703, 
    -233.333282470703, 
    -205.595306396484, 
    -125.054748535156, 
    -154.885864257812, 
    -159.750381469727, 
    -231.393081665039, 
    -665.491333007812, 
    -427.586334228516, 
    262.285797119141, 
    8.1501350402832, 
    516.9111328125, 
    80.4749984741211, 
    674.777770996094, 
    735.972229003906, 
    669.002807617188, 
    126.216178894043, 
    -26.5987014770508, 
    670.274108886719, 
    354.052764892578, 
    463.586120605469, 
    687.347229003906, 
    922.099975585938, 
    620.391662597656, 
    444.477783203125, 
    -269.986022949219, 
    -459.969207763672, 
    -342.547210693359, 
    -201.759750366211, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -203.549819946289, 
    -248.333221435547, 
    -200, 
    -200, 
    -200, 
    -200, 
    -204.042755126953, 
    -200, 
    -200, 
    -200,
  
    -3424.79956054688, 
    -3404.33544921875, 
    -3392.96728515625, 
    -3381.38940429688, 
    -3354.701171875, 
    -3328.88159179688, 
    -3225.798828125, 
    -3132.54028320312, 
    -3070.05541992188, 
    -3020.14575195312, 
    -2981.98852539062, 
    -2974.42724609375, 
    -2934.70336914062, 
    -2913.09106445312, 
    -2905.5029296875, 
    -2824.17529296875, 
    -2724.78857421875, 
    -2617.02612304688, 
    -2508.80688476562, 
    -2313.29516601562, 
    -1749.95336914062, 
    -805.136474609375, 
    -417.282287597656, 
    -112.803977966309, 
    -352.990997314453, 
    -92.727165222168, 
    -55.5559768676758, 
    -83.5053558349609, 
    -321.870697021484, 
    -166.47102355957, 
    -102.255279541016, 
    -88.6652984619141, 
    -95.9203567504883, 
    -146.673309326172, 
    -259.228088378906, 
    -235.484512329102, 
    -142.422439575195, 
    -210.819534301758, 
    -155.337188720703, 
    -17.765625, 
    24.4268531799316, 
    74.5357666015625, 
    114.431686401367, 
    168.634887695312, 
    165.898788452148, 
    -59.1920394897461, 
    -269.422576904297, 
    -110.072364807129, 
    -85.1538238525391, 
    -54.9331130981445, 
    -49.6671409606934, 
    -31.0796432495117, 
    -30.1196384429932, 
    -24.9892234802246, 
    -35.3791007995605, 
    -193.058700561523, 
    -454.213684082031, 
    -344.710113525391, 
    -229.679870605469, 
    -143.132293701172, 
    -144.759323120117, 
    -185.607299804688, 
    -225.625228881836, 
    -197.973098754883, 
    -146.870803833008, 
    -154.31379699707, 
    -176.566390991211, 
    -255.802429199219, 
    -320.149261474609, 
    -485.828521728516, 
    -506.675720214844, 
    -348.545196533203, 
    -302.353637695312, 
    -255.821533203125, 
    -276.087249755859, 
    -279.381927490234, 
    -303.722137451172, 
    -315.645965576172, 
    -335.283142089844, 
    -307.918853759766, 
    -286.0693359375, 
    -396.243072509766, 
    -613.005249023438, 
    -615.842041015625, 
    -356.519104003906, 
    -303.373687744141, 
    -361.273986816406, 
    -438.689117431641, 
    -522.258850097656, 
    -551.789794921875, 
    -625.845092773438, 
    -634.4091796875, 
    -623.49072265625, 
    -368.362762451172, 
    -369.700500488281, 
    -207.191635131836, 
    -135.632888793945, 
    -169.677871704102, 
    -204.51123046875, 
    -568.435546875, 
    -716.079833984375, 
    -437.837188720703, 
    62.5857582092285, 
    431.922210693359, 
    624.141662597656, 
    672.899963378906, 
    728.174987792969, 
    757.16943359375, 
    546.808349609375, 
    661.825012207031, 
    -542.026062011719, 
    588.375, 
    392.050018310547, 
    648.097229003906, 
    521.377807617188, 
    801.200012207031, 
    459.997222900391, 
    345.625, 
    -282.534515380859, 
    -303.628784179688, 
    -244.540542602539, 
    -217.74397277832, 
    -207.445663452148, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -204.030014038086, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3406.84716796875, 
    -3384.2509765625, 
    -3364.02001953125, 
    -3353.70581054688, 
    -3338.1005859375, 
    -3266.2607421875, 
    -3179.75146484375, 
    -3061.384765625, 
    -2995.02685546875, 
    -2949.16650390625, 
    -2920.65576171875, 
    -2941.26806640625, 
    -2895.15600585938, 
    -2844.66137695312, 
    -2807.42309570312, 
    -1914.78283691406, 
    -1042.77758789062, 
    -1397.02380371094, 
    -1862.607421875, 
    -1323.03833007812, 
    -1155.44958496094, 
    -238.581985473633, 
    -149.334671020508, 
    -76.7854690551758, 
    -331.624450683594, 
    -211.298736572266, 
    -123.199844360352, 
    -98.9047088623047, 
    -78.991584777832, 
    -32.6680793762207, 
    -28.2192535400391, 
    31.748140335083, 
    47.5167579650879, 
    4.1147985458374, 
    -65.4544906616211, 
    -65.4117584228516, 
    38.7180061340332, 
    17.7728748321533, 
    -6.86234903335571, 
    218.919372558594, 
    472.683013916016, 
    219.96110534668, 
    683.469421386719, 
    657.480590820312, 
    710.430541992188, 
    85.5687026977539, 
    -10.3989906311035, 
    54.3343734741211, 
    182.574996948242, 
    50.8456230163574, 
    -55.3117523193359, 
    -44.3923301696777, 
    -41.5593795776367, 
    -69.5706329345703, 
    -178.781234741211, 
    -259.811248779297, 
    -299.011077880859, 
    -308.416870117188, 
    -240.183044433594, 
    -202.297805786133, 
    -181.84098815918, 
    -207.332946777344, 
    -251.58447265625, 
    -136.201202392578, 
    -103.978004455566, 
    -123.661796569824, 
    -113.645561218262, 
    -185.094451904297, 
    -275.653198242188, 
    -512.633850097656, 
    -537.376037597656, 
    -375.379577636719, 
    -291.765716552734, 
    -227.319046020508, 
    -237.651885986328, 
    -231.921615600586, 
    -240.923049926758, 
    -245.077453613281, 
    -302.525848388672, 
    -267.745880126953, 
    -195.343399047852, 
    -209.720718383789, 
    -480.440612792969, 
    -713.800903320312, 
    -445.529052734375, 
    -258.929779052734, 
    -309.528564453125, 
    -379.263458251953, 
    -522.845764160156, 
    -599.911804199219, 
    -651.731689453125, 
    -684.265930175781, 
    -740.092163085938, 
    -604.115417480469, 
    -554.810363769531, 
    -527.481384277344, 
    -359.878570556641, 
    -304.358215332031, 
    -384.551910400391, 
    -408.327972412109, 
    -616.888610839844, 
    -42.7857475280762, 
    64.622184753418, 
    434.316650390625, 
    797.658325195312, 
    936.163879394531, 
    619.599975585938, 
    480.491668701172, 
    471.952789306641, 
    84.4269485473633, 
    -230.191680908203, 
    700.79443359375, 
    888.488891601562, 
    710.561096191406, 
    705.144409179688, 
    613.161071777344, 
    521.497253417969, 
    398.644439697266, 
    -221.566757202148, 
    -281.864379882812, 
    -201.395065307617, 
    -201.836090087891, 
    -240.130081176758, 
    -200, 
    -200, 
    -243.578506469727, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -201.292526245117, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3373.57934570312, 
    -3327.28295898438, 
    -3342.71997070312, 
    -3333.50268554688, 
    -3299.25366210938, 
    -3198.88452148438, 
    -3096.87377929688, 
    -3006.587890625, 
    -2944.82861328125, 
    -2893.74365234375, 
    -2862.41748046875, 
    -2868.82250976562, 
    -2789.8818359375, 
    -2570.076171875, 
    -1112.57678222656, 
    -184.974746704102, 
    -112.08854675293, 
    -112.865020751953, 
    -329.331146240234, 
    -114.582458496094, 
    -248.165634155273, 
    -184.109146118164, 
    -171.754776000977, 
    -101.598709106445, 
    -68.0327835083008, 
    12.8871555328369, 
    0.317923009395599, 
    65.1972198486328, 
    169.530548095703, 
    78.9148788452148, 
    168.734527587891, 
    171.384368896484, 
    139.057678222656, 
    186.077774047852, 
    217.522216796875, 
    103.016662597656, 
    345.341674804688, 
    365.041656494141, 
    386.394439697266, 
    530.386108398438, 
    1155.14440917969, 
    647.597229003906, 
    1102.77770996094, 
    622.538879394531, 
    1231.57775878906, 
    586.327758789062, 
    197.297973632812, 
    307.294860839844, 
    438.130554199219, 
    500.274993896484, 
    293.324981689453, 
    69.2773361206055, 
    9.09448337554932, 
    -51.4614410400391, 
    -200.093200683594, 
    -395.575805664062, 
    -528.962585449219, 
    -293.885620117188, 
    -195.084915161133, 
    -167.758911132812, 
    -146.371719360352, 
    -236.751937866211, 
    -143.214553833008, 
    -83.0682678222656, 
    -83.216911315918, 
    -83.9175872802734, 
    -82.1017532348633, 
    -94.1505508422852, 
    -155.793273925781, 
    -519.860046386719, 
    -552.059631347656, 
    -356.160186767578, 
    -244.996047973633, 
    -188.451507568359, 
    -195.524490356445, 
    -198.031539916992, 
    -198.97624206543, 
    -281.121002197266, 
    -291.284240722656, 
    -237.317276000977, 
    -179.288803100586, 
    -145.74137878418, 
    -273.520111083984, 
    -782.205383300781, 
    -586.868774414062, 
    -218.490325927734, 
    -183.228179931641, 
    -277.538635253906, 
    -471.287872314453, 
    -615.658996582031, 
    -696.23193359375, 
    -754.962219238281, 
    -747.490539550781, 
    -777.593322753906, 
    -801.099670410156, 
    -836.225830078125, 
    -970.42919921875, 
    -994.220031738281, 
    -821.658203125, 
    -580.005065917969, 
    -463.271484375, 
    -79.2942428588867, 
    140.025054931641, 
    732.111083984375, 
    900.20556640625, 
    609.441650390625, 
    589.763854980469, 
    513.186096191406, 
    496.700012207031, 
    392.700134277344, 
    65.7832565307617, 
    567.252807617188, 
    803.983337402344, 
    689.799987792969, 
    742.369445800781, 
    654.766662597656, 
    412.091674804688, 
    252.341659545898, 
    -217.627151489258, 
    -318.314575195312, 
    -192.97900390625, 
    -200.206802368164, 
    -234.554336547852, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3323.328125, 
    -3280.41967773438, 
    -3279.00903320312, 
    -3299.50244140625, 
    -3237.09301757812, 
    -3127.67236328125, 
    -3046.484375, 
    -2938.34057617188, 
    -2866.99438476562, 
    -2821.06909179688, 
    -2752.93676757812, 
    -2627.26782226562, 
    -2415.25439453125, 
    -990.977783203125, 
    -218.997833251953, 
    -180.016006469727, 
    -180.474807739258, 
    -146.304702758789, 
    -179.330780029297, 
    -115.654945373535, 
    -70.9109649658203, 
    -44.6721305847168, 
    9.43384838104248, 
    -15.1339511871338, 
    15.4294548034668, 
    244.975006103516, 
    242.505554199219, 
    612.75, 
    563.511108398438, 
    440.613891601562, 
    528.355590820312, 
    321.763885498047, 
    330.654846191406, 
    35.6410255432129, 
    198.969436645508, 
    132.432144165039, 
    392.299987792969, 
    550.466674804688, 
    557.547241210938, 
    399.311126708984, 
    963.408325195312, 
    686.897216796875, 
    1423.5, 
    1569.73889160156, 
    632.430541992188, 
    375.555541992188, 
    210.261108398438, 
    750.197204589844, 
    882.738891601562, 
    717.775024414062, 
    404.29443359375, 
    115.516662597656, 
    113.64722442627, 
    56.9269943237305, 
    0.368709057569504, 
    -76.266845703125, 
    -346.805603027344, 
    -767.0029296875, 
    -203.799591064453, 
    -113.951728820801, 
    -196.60888671875, 
    -57.5709762573242, 
    225.001922607422, 
    216.871673583984, 
    193.02555847168, 
    -84.8679885864258, 
    -151.702438354492, 
    -109.727615356445, 
    -316.739807128906, 
    -484.685943603516, 
    -532.69775390625, 
    -326.317230224609, 
    -198.541213989258, 
    -207.935775756836, 
    -186.786209106445, 
    -152.265441894531, 
    -195.229721069336, 
    -246.934997558594, 
    -320.226135253906, 
    -192.007217407227, 
    -206.371704101562, 
    -139.971420288086, 
    -327.187286376953, 
    -749.946228027344, 
    -824.060974121094, 
    -540.552673339844, 
    -234.236557006836, 
    -127.442993164062, 
    -210.651062011719, 
    -536.307067871094, 
    -764.184509277344, 
    -788.632751464844, 
    -814.956176757812, 
    -776.016479492188, 
    -793.405700683594, 
    -813.432067871094, 
    -770.638610839844, 
    -494.005676269531, 
    -432.259429931641, 
    -217.759963989258, 
    -32.7070693969727, 
    2.27411460876465, 
    369.236114501953, 
    927.819458007812, 
    754.174987792969, 
    704.113891601562, 
    632.983337402344, 
    481.322235107422, 
    448.211120605469, 
    112.944442749023, 
    224.683334350586, 
    619.305541992188, 
    735.0361328125, 
    665.652770996094, 
    663.049987792969, 
    621.258361816406, 
    526.744445800781, 
    286.475006103516, 
    83.22265625, 
    -281.086761474609, 
    -189.556365966797, 
    -192.675109863281, 
    -216.131637573242, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3291.16186523438, 
    -3272.29956054688, 
    -3243.64990234375, 
    -3252.42578125, 
    -3172.818359375, 
    -3053.95385742188, 
    -2946.59375, 
    -2937.95361328125, 
    -2808.71899414062, 
    -2685.38330078125, 
    -1740.6748046875, 
    -216.447463989258, 
    -180.805313110352, 
    -186.657852172852, 
    -113.125175476074, 
    -102.454330444336, 
    -91.8999710083008, 
    -39.1476554870605, 
    -23.4191188812256, 
    0.738058149814606, 
    183.141662597656, 
    300.70556640625, 
    151.002777099609, 
    310.377777099609, 
    465.161102294922, 
    488.325012207031, 
    825.497192382812, 
    999.055541992188, 
    1152.29724121094, 
    673.761108398438, 
    784.308837890625, 
    736.5361328125, 
    407.373107910156, 
    67.0569839477539, 
    296.597229003906, 
    570.011108398438, 
    323.549987792969, 
    639.227783203125, 
    570.822204589844, 
    585.49169921875, 
    611.788879394531, 
    951.733337402344, 
    1522.52502441406, 
    1261.57775878906, 
    527.174987792969, 
    387.088897705078, 
    439.005554199219, 
    463.908355712891, 
    1044.73889160156, 
    447.16943359375, 
    330.658325195312, 
    177.987197875977, 
    257.513885498047, 
    126.25, 
    22.8920955657959, 
    69.4306488037109, 
    -66.6232681274414, 
    -364.366668701172, 
    -608.412902832031, 
    -305.443908691406, 
    308.904327392578, 
    116.792915344238, 
    429.149993896484, 
    704.680541992188, 
    647.344421386719, 
    737.122192382812, 
    -110.855628967285, 
    -211.4775390625, 
    -381.073760986328, 
    -535.269836425781, 
    -481.38671875, 
    -274.040588378906, 
    -100.470252990723, 
    2.91175580024719, 
    197.88330078125, 
    -103.770149230957, 
    -165.675247192383, 
    -191.490905761719, 
    -287.687713623047, 
    -260.181518554688, 
    -201.141998291016, 
    -282.81884765625, 
    -447.413909912109, 
    -512.576354980469, 
    -609.584106445312, 
    -811.715026855469, 
    -603.717895507812, 
    -322.168701171875, 
    -334.610443115234, 
    -341.512725830078, 
    -824.57275390625, 
    -742.340881347656, 
    -741.998046875, 
    -431.623077392578, 
    -447.952453613281, 
    -296.987579345703, 
    -217.753768920898, 
    -197.514511108398, 
    -146.0419921875, 
    -40.1305389404297, 
    16.1736736297607, 
    207.891662597656, 
    726.494445800781, 
    547.4111328125, 
    584.936096191406, 
    684.380554199219, 
    564.033325195312, 
    617.991638183594, 
    479.386108398438, 
    541.302734375, 
    572.277770996094, 
    645.755554199219, 
    713.933349609375, 
    648.91943359375, 
    615.633361816406, 
    421.963897705078, 
    426, 
    266.674987792969, 
    62.6994743347168, 
    -301.420501708984, 
    -173.60466003418, 
    -165.022079467773, 
    -200.271270751953, 
    -206.075637817383, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -294.40673828125,
  
    -3247.01733398438, 
    -3201.66357421875, 
    -3172.455078125, 
    -3178.95654296875, 
    -3150.4794921875, 
    -2987.37084960938, 
    -2849.1640625, 
    -2795.40405273438, 
    -2473.1845703125, 
    -819.623840332031, 
    -150.079147338867, 
    -178.637145996094, 
    -178.829803466797, 
    -99.9018783569336, 
    -88.9048919677734, 
    0.972452640533447, 
    134.030380249023, 
    100.805557250977, 
    205.543518066406, 
    289.697235107422, 
    476.022216796875, 
    742.255554199219, 
    816.3388671875, 
    698.841674804688, 
    1061.13061523438, 
    695.802795410156, 
    698.861083984375, 
    1149.19165039062, 
    799.313842773438, 
    548.569458007812, 
    642.322204589844, 
    376.108337402344, 
    760.50830078125, 
    308.29443359375, 
    218.53889465332, 
    243.400009155273, 
    344.575012207031, 
    607.219421386719, 
    589.827758789062, 
    790.127746582031, 
    951.702758789062, 
    1590.41662597656, 
    975.575012207031, 
    909.966674804688, 
    567.138854980469, 
    177.980087280273, 
    374.674987792969, 
    679.322204589844, 
    819.325012207031, 
    281.594451904297, 
    439.130554199219, 
    159.941619873047, 
    128.769439697266, 
    130.66667175293, 
    54.0873680114746, 
    74.478874206543, 
    59.6068992614746, 
    -290.285217285156, 
    -287.237976074219, 
    -453.625732421875, 
    409.056823730469, 
    635.075012207031, 
    640.238891601562, 
    1190.69165039062, 
    1082.00549316406, 
    521.977783203125, 
    -289.916290283203, 
    79.6393051147461, 
    496.473175048828, 
    -578.41064453125, 
    -464.017578125, 
    -140.333770751953, 
    65.7457580566406, 
    465.058349609375, 
    390.166687011719, 
    88.3228302001953, 
    -42.5026550292969, 
    -70.5343399047852, 
    -253.789260864258, 
    -171.38053894043, 
    -140.397308349609, 
    -54.1913528442383, 
    -241.53874206543, 
    -114.423622131348, 
    -149.691268920898, 
    -125.247177124023, 
    -231.297592163086, 
    -181.842315673828, 
    -161.060668945312, 
    -224.7568359375, 
    -135.714294433594, 
    -166.635971069336, 
    -238.981201171875, 
    -231.353042602539, 
    -239.563232421875, 
    -188.017761230469, 
    -198.937301635742, 
    -188.275436401367, 
    -16.5351123809814, 
    29.3990440368652, 
    547.502319335938, 
    148.625, 
    385.636108398438, 
    667.947204589844, 
    548.847229003906, 
    589.122253417969, 
    600.252746582031, 
    582.6611328125, 
    574.936096191406, 
    548.966674804688, 
    685.038879394531, 
    584.991638183594, 
    623.083312988281, 
    544.591674804688, 
    482.833312988281, 
    378.258331298828, 
    202.925003051758, 
    242.088882446289, 
    -66.8208770751953, 
    -321.316619873047, 
    -166.642974853516, 
    -124.384796142578, 
    -181.676727294922, 
    -234.062026977539, 
    -201.894409179688, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3165.8916015625, 
    -3138.28344726562, 
    -3143.4482421875, 
    -2998.39770507812, 
    -3019.89624023438, 
    -3006.35693359375, 
    -2808.65356445312, 
    -2626.42749023438, 
    -459.353851318359, 
    -197.335693359375, 
    -157.37939453125, 
    -152.135375976562, 
    -97.4483032226562, 
    -30.6621017456055, 
    244.869445800781, 
    300.075012207031, 
    502.019439697266, 
    423.929870605469, 
    444.777801513672, 
    754.33056640625, 
    804.513854980469, 
    1090.73889160156, 
    1125.63049316406, 
    1207.06115722656, 
    1180.26391601562, 
    832.836120605469, 
    784.166687011719, 
    988.058349609375, 
    920.608337402344, 
    520.994445800781, 
    553.04443359375, 
    635.791687011719, 
    306.280456542969, 
    393.401947021484, 
    715.333312988281, 
    899.677795410156, 
    619.622192382812, 
    623.822204589844, 
    568.219421386719, 
    306.441650390625, 
    1058.43603515625, 
    1235.56665039062, 
    1214.81945800781, 
    1022.51940917969, 
    598.052795410156, 
    504.338897705078, 
    317.530578613281, 
    431.094451904297, 
    486.647216796875, 
    506.119445800781, 
    178.908157348633, 
    368.211120605469, 
    164.58610534668, 
    146.680557250977, 
    159.661117553711, 
    261.25, 
    59.2524337768555, 
    -225.39778137207, 
    -337.124145507812, 
    -499.863372802734, 
    39.7258224487305, 
    1037.79724121094, 
    1155.34997558594, 
    1195.02221679688, 
    1342.64440917969, 
    96.2559432983398, 
    673.55712890625, 
    1108.23608398438, 
    351.090179443359, 
    -684.2919921875, 
    -306.240234375, 
    -197.297286987305, 
    456.480560302734, 
    354.558349609375, 
    625.255554199219, 
    338.841674804688, 
    730.069458007812, 
    187.83821105957, 
    368.861114501953, 
    341.594451904297, 
    59.7456550598145, 
    0.703871309757233, 
    45.8743705749512, 
    34.1866722106934, 
    9.81857204437256, 
    37.4093475341797, 
    60.3064842224121, 
    -19.2907085418701, 
    -47.9601440429688, 
    -32.8664970397949, 
    -37.1750717163086, 
    -3.71728897094727, 
    -23.1862640380859, 
    -104.131278991699, 
    -112.148475646973, 
    -143.943771362305, 
    -81.1474990844727, 
    35.2549057006836, 
    164.441360473633, 
    176.483337402344, 
    302.911102294922, 
    275.269439697266, 
    344.416656494141, 
    619.799987792969, 
    570.269409179688, 
    553.686096191406, 
    535.961120605469, 
    525.694458007812, 
    571.611145019531, 
    593.230529785156, 
    642.194458007812, 
    609.563903808594, 
    611.358337402344, 
    568.383361816406, 
    521.030578613281, 
    490.991668701172, 
    395.969451904297, 
    111.917663574219, 
    -179.356170654297, 
    -344.709014892578, 
    -182.231018066406, 
    -97.2828216552734, 
    -183.083648681641, 
    -236.857543945312, 
    -269.237152099609, 
    -233.812484741211, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -3099.91723632812, 
    -2999.57104492188, 
    -3069.333984375, 
    -2985.2724609375, 
    -2908.78979492188, 
    -2824.80395507812, 
    -2777.78344726562, 
    -792.797912597656, 
    -129.661392211914, 
    -104.372703552246, 
    14.595401763916, 
    11.7658395767212, 
    285.387939453125, 
    267.636108398438, 
    556.441650390625, 
    486.113891601562, 
    846.3388671875, 
    522.113891601562, 
    996.755554199219, 
    1060.29724121094, 
    1095.74438476562, 
    1225.88061523438, 
    1317.79443359375, 
    1398.68334960938, 
    1473.11669921875, 
    1362.5888671875, 
    1166.44165039062, 
    1122.12780761719, 
    894.694458007812, 
    796.502746582031, 
    564.741638183594, 
    514.744445800781, 
    800.125, 
    863.577758789062, 
    907.283325195312, 
    896.094421386719, 
    834.427734375, 
    803.297241210938, 
    625, 
    664.133361816406, 
    1002.52502441406, 
    1268.19165039062, 
    1105.83605957031, 
    957.352783203125, 
    782.247253417969, 
    348.113891601562, 
    191.619445800781, 
    299.261108398438, 
    514.019470214844, 
    412.41943359375, 
    97.5772399902344, 
    76.0052947998047, 
    245.941665649414, 
    22.5887603759766, 
    137.819595336914, 
    22.4038600921631, 
    -152.294616699219, 
    -106.580528259277, 
    -346.723022460938, 
    -379.569732666016, 
    -199.436172485352, 
    467.397216796875, 
    522.241638183594, 
    -50.1182403564453, 
    -458.946533203125, 
    51.3830642700195, 
    361.911102294922, 
    1042.71105957031, 
    -366.237915039062, 
    -641.374206542969, 
    454.941955566406, 
    -151.168853759766, 
    20.9619579315186, 
    89.1762924194336, 
    798.74169921875, 
    1047.9638671875, 
    570.200012207031, 
    348.977783203125, 
    181.022216796875, 
    168.952774047852, 
    -3.69295287132263, 
    226.816665649414, 
    25.0646228790283, 
    52.0526809692383, 
    72.5890960693359, 
    52.2329292297363, 
    48.4499702453613, 
    27.4410190582275, 
    38.3849868774414, 
    64.8364715576172, 
    60.8108749389648, 
    -1.94466364383698, 
    89.5976638793945, 
    -353.733337402344, 
    73.0694427490234, 
    230.612030029297, 
    114.754295349121, 
    108.177780151367, 
    217.127777099609, 
    265.497222900391, 
    370.497222900391, 
    268.716674804688, 
    306.813873291016, 
    348.819427490234, 
    509.705535888672, 
    550.963928222656, 
    559.211120605469, 
    541.433349609375, 
    560.002807617188, 
    551.477783203125, 
    564.322204589844, 
    586.533325195312, 
    546.772216796875, 
    509.072235107422, 
    478.811126708984, 
    389.247222900391, 
    264.133331298828, 
    12.5861110687256, 
    -115.136367797852, 
    -297.219207763672, 
    -184.536560058594, 
    -94.7271499633789, 
    -104.862686157227, 
    -244.293762207031, 
    -340.797149658203, 
    -296.457397460938, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -2876.41870117188, 
    -2948.89697265625, 
    -2918.60107421875, 
    -2892.61791992188, 
    -2821.91479492188, 
    -2725.8515625, 
    -2058.83813476562, 
    -177.57145690918, 
    -122.362129211426, 
    -71.5562973022461, 
    60.888744354248, 
    14.5082845687866, 
    452.286102294922, 
    426.675018310547, 
    733.163879394531, 
    684.566650390625, 
    1020.95001220703, 
    884.524963378906, 
    1064.59167480469, 
    1106.27783203125, 
    1262.37780761719, 
    1399.66662597656, 
    1479.92224121094, 
    1360.21948242188, 
    1377.7138671875, 
    1239.0166015625, 
    1043.73889160156, 
    768.911071777344, 
    629.41943359375, 
    458.383331298828, 
    772.297241210938, 
    1017.65551757812, 
    986.79443359375, 
    896.755554199219, 
    1045.77221679688, 
    1001.51666259766, 
    810.194458007812, 
    756.825012207031, 
    719.163879394531, 
    701.24169921875, 
    780.630554199219, 
    898.694458007812, 
    1009.83337402344, 
    813.908325195312, 
    490.486114501953, 
    287.741668701172, 
    292.458343505859, 
    324.297210693359, 
    465.827758789062, 
    206.544448852539, 
    362.891662597656, 
    204.786117553711, 
    54.6957550048828, 
    262.691680908203, 
    121.51782989502, 
    27.0976734161377, 
    -212.821472167969, 
    -285.021942138672, 
    -331.740478515625, 
    -329.559234619141, 
    -250.595458984375, 
    50.9881973266602, 
    124.750305175781, 
    -364.750335693359, 
    533.552795410156, 
    724.138916015625, 
    1058.59997558594, 
    1050.87561035156, 
    -522.01513671875, 
    -538.286254882812, 
    213.42707824707, 
    -144.402481079102, 
    -10.5305671691895, 
    -181.972579956055, 
    890.686096191406, 
    897.647216796875, 
    890.550048828125, 
    452.347229003906, 
    647.077758789062, 
    202.938888549805, 
    -19.7375144958496, 
    364.836120605469, 
    304.33056640625, 
    245.730545043945, 
    333.263885498047, 
    234.747222900391, 
    312.316680908203, 
    363.680572509766, 
    92.6555557250977, 
    162.31266784668, 
    130.099990844727, 
    203.441665649414, 
    56.0444450378418, 
    42.4194450378418, 
    151.761108398438, 
    366.908325195312, 
    63.7805557250977, 
    264.308319091797, 
    150.327774047852, 
    354.188873291016, 
    284.54443359375, 
    297.852783203125, 
    398.399993896484, 
    359.269439697266, 
    454.655548095703, 
    392.238891601562, 
    422.625, 
    408.108337402344, 
    372.377777099609, 
    320.899993896484, 
    431.658325195312, 
    506.966674804688, 
    490.988891601562, 
    438.922210693359, 
    372.491668701172, 
    321.602783203125, 
    224.741668701172, 
    27.9972229003906, 
    -115.880554199219, 
    -236.2314453125, 
    -199.759902954102, 
    -117.483512878418, 
    43.3142967224121, 
    227.458343505859, 
    -194.045349121094, 
    -354.394958496094, 
    -205.787536621094, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -2784.884765625, 
    -2807.42553710938, 
    -2643.05883789062, 
    -2614.61450195312, 
    -2689.24682617188, 
    -2014.10913085938, 
    -487.392547607422, 
    -116.244445800781, 
    -151.229965209961, 
    -70.9679870605469, 
    44.8278121948242, 
    176.763885498047, 
    642.099975585938, 
    983.083312988281, 
    1139.94165039062, 
    1020.18609619141, 
    1092.08325195312, 
    1060.26940917969, 
    985.2138671875, 
    1093.48889160156, 
    1210.96948242188, 
    1499.34167480469, 
    1339.89440917969, 
    1202.09997558594, 
    1161.08056640625, 
    858.533325195312, 
    1157.79162597656, 
    899.791687011719, 
    720.694458007812, 
    846.105590820312, 
    790.788879394531, 
    1040.94165039062, 
    961.422241210938, 
    797.769470214844, 
    793.08056640625, 
    758.880554199219, 
    654.4638671875, 
    646.477783203125, 
    584.472229003906, 
    519.902770996094, 
    559.450012207031, 
    743.647216796875, 
    895.325012207031, 
    742.316650390625, 
    449.936096191406, 
    437.383331298828, 
    265.380554199219, 
    403.399993896484, 
    561.358337402344, 
    401.894439697266, 
    267.247222900391, 
    185.850006103516, 
    240.925003051758, 
    215.130554199219, 
    313.672210693359, 
    235.513885498047, 
    220.762985229492, 
    219.739837646484, 
    -153.390991210938, 
    -356.227325439453, 
    -244.714477539062, 
    -264.556762695312, 
    -491.404937744141, 
    125.025810241699, 
    879.513916015625, 
    882.549987792969, 
    653.423278808594, 
    -340.41796875, 
    -203.129379272461, 
    -357.649169921875, 
    341.233245849609, 
    596.324096679688, 
    -259.041625976562, 
    1233.73889160156, 
    686.143859863281, 
    1032.72778320312, 
    1418.7861328125, 
    842.072204589844, 
    609.047241210938, 
    199.411117553711, 
    223.508331298828, 
    266.269439697266, 
    311.938903808594, 
    231.824996948242, 
    238.397216796875, 
    302.691680908203, 
    282.708312988281, 
    81.4805526733398, 
    244.002777099609, 
    221.397216796875, 
    166.169448852539, 
    195.08610534668, 
    53.8583335876465, 
    252.074996948242, 
    196.544448852539, 
    355.574981689453, 
    426.791656494141, 
    228.952774047852, 
    276.388885498047, 
    276.416656494141, 
    159.152770996094, 
    255.697219848633, 
    468.486114501953, 
    405.930572509766, 
    317.497222900391, 
    245.652786254883, 
    192.20832824707, 
    204.883331298828, 
    236.511108398438, 
    363.019439697266, 
    439.616668701172, 
    446.105560302734, 
    435.316680908203, 
    347.111114501953, 
    289.991668701172, 
    234.399993896484, 
    125.633331298828, 
    12.0083332061768, 
    -138.897216796875, 
    -178.608337402344, 
    -79.5645141601562, 
    -46.7414016723633, 
    468.302795410156, 
    503.761108398438, 
    326.652770996094, 
    -250.320816040039, 
    -330.609588623047, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -337.667724609375, 
    -327.206146240234,
  
    -2563.91015625, 
    -2275.16455078125, 
    -2252.02197265625, 
    -2080.02465820312, 
    -2339.001953125, 
    -1933.97998046875, 
    -324.292175292969, 
    -343.000244140625, 
    -444.420104980469, 
    -41.2129249572754, 
    10.7336254119873, 
    361.583343505859, 
    1078.35559082031, 
    1284.0166015625, 
    1339.95275878906, 
    1201.22778320312, 
    1052.0166015625, 
    893.336120605469, 
    719.450012207031, 
    863.724975585938, 
    1222.50549316406, 
    1219.63330078125, 
    1170.18054199219, 
    947.647216796875, 
    1001.24719238281, 
    964.266662597656, 
    1015.63055419922, 
    880.377746582031, 
    612.408325195312, 
    508.858337402344, 
    612.138916015625, 
    840.988891601562, 
    816.041687011719, 
    625.7861328125, 
    560.474975585938, 
    576.622192382812, 
    491.433349609375, 
    570.344421386719, 
    564.224975585938, 
    583.530578613281, 
    611.172241210938, 
    713.652770996094, 
    724.7861328125, 
    656.647216796875, 
    556.113891601562, 
    397.949981689453, 
    218.180557250977, 
    359.047210693359, 
    575.95556640625, 
    517.70556640625, 
    398.825012207031, 
    415.922210693359, 
    429.580535888672, 
    329.963897705078, 
    347.997222900391, 
    317.799987792969, 
    229.686111450195, 
    69.6333312988281, 
    -378.818542480469, 
    437.008331298828, 
    97.5261611938477, 
    -1.74831306934357, 
    164.120147705078, 
    151.862991333008, 
    917.069458007812, 
    576.180297851562, 
    -182.76708984375, 
    -497.961303710938, 
    56.2521934509277, 
    -314.82080078125, 
    359.518371582031, 
    1205.70178222656, 
    336.268951416016, 
    792.174987792969, 
    1391.53051757812, 
    1037.68334960938, 
    1829.6611328125, 
    1199.43334960938, 
    772.672241210938, 
    415.038879394531, 
    465.063903808594, 
    400.969451904297, 
    265.063873291016, 
    205.361114501953, 
    28.2972221374512, 
    138.572219848633, 
    145.938888549805, 
    164.66667175293, 
    365.288879394531, 
    327.608337402344, 
    256.450012207031, 
    229.222229003906, 
    254.330551147461, 
    278.286102294922, 
    228.25, 
    361.466674804688, 
    447.161102294922, 
    340.54443359375, 
    321.561126708984, 
    333.172210693359, 
    357.211120605469, 
    203.183334350586, 
    340.344451904297, 
    316.163879394531, 
    245.925003051758, 
    200.266677856445, 
    100.166664123535, 
    156.730560302734, 
    422.230560302734, 
    456.661102294922, 
    369.405548095703, 
    324.877777099609, 
    299.341674804688, 
    253.33610534668, 
    221.766662597656, 
    178.83610534668, 
    57.1111106872559, 
    -78.3111114501953, 
    -101.888885498047, 
    -281.841674804688, 
    -35.1777801513672, 
    330.466979980469, 
    516.447204589844, 
    422.263885498047, 
    485.911102294922, 
    -135.188217163086, 
    -374.437225341797, 
    -200, 
    -200, 
    -209.727310180664, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -2435.04809570312, 
    -2157.24829101562, 
    -2084.64721679688, 
    -1594.3525390625, 
    -1358.76721191406, 
    -452.794006347656, 
    -149.643936157227, 
    -481.958984375, 
    -91.1504211425781, 
    1.47775566577911, 
    230.894439697266, 
    552.522216796875, 
    1123.8583984375, 
    1249.46667480469, 
    1271.56665039062, 
    1162.94445800781, 
    857.291687011719, 
    742.494445800781, 
    688.036071777344, 
    812.247192382812, 
    1182.69995117188, 
    1272.125, 
    1044.91943359375, 
    982.813903808594, 
    972.447204589844, 
    971.730529785156, 
    875.433349609375, 
    758.147216796875, 
    522.322204589844, 
    484.611114501953, 
    673.072204589844, 
    814.777770996094, 
    853.799987792969, 
    898.991638183594, 
    732.6611328125, 
    549.761108398438, 
    574.702758789062, 
    580.99169921875, 
    492.541656494141, 
    493.016662597656, 
    511.572204589844, 
    613.70556640625, 
    712.508361816406, 
    639.04443359375, 
    424.308349609375, 
    299.780548095703, 
    177.202774047852, 
    278.522216796875, 
    497.344451904297, 
    513.613891601562, 
    505.649993896484, 
    410.838897705078, 
    399.238891601562, 
    262.094451904297, 
    18.1249980926514, 
    115.655555725098, 
    176.871627807617, 
    293.737396240234, 
    -291.79248046875, 
    -176.753204345703, 
    304.466369628906, 
    255.540435791016, 
    118.599433898926, 
    184.422225952148, 
    645.505554199219, 
    170.38264465332, 
    37.8079490661621, 
    -53.3477973937988, 
    498.942016601562, 
    365.333343505859, 
    652.172241210938, 
    186.048828125, 
    757.045715332031, 
    1693.53051757812, 
    1508.90551757812, 
    1849.74450683594, 
    1219.67224121094, 
    1192.69165039062, 
    693.936096191406, 
    491.658325195312, 
    364.072235107422, 
    378.5, 
    366.313873291016, 
    375.869445800781, 
    267.25, 
    200.697219848633, 
    160.811111450195, 
    145.022216796875, 
    172.988891601562, 
    256.95556640625, 
    188.716674804688, 
    325.944458007812, 
    416.330535888672, 
    403.5888671875, 
    364.625, 
    516.422180175781, 
    633, 
    518.888916015625, 
    501.844421386719, 
    237.716659545898, 
    300.366668701172, 
    186.255554199219, 
    179.719451904297, 
    129.638885498047, 
    179.930557250977, 
    81.0138931274414, 
    135.027770996094, 
    308.311126708984, 
    371.788879394531, 
    296.225006103516, 
    147.122222900391, 
    170.544448852539, 
    182.411117553711, 
    130.858337402344, 
    137.269439697266, 
    93.533332824707, 
    45.2333335876465, 
    -25.8861103057861, 
    -67.0500030517578, 
    -108.52222442627, 
    337.255554199219, 
    397.572235107422, 
    466.997222900391, 
    657.052795410156, 
    724.166687011719, 
    257.387786865234, 
    -334.297241210938, 
    -307.228363037109, 
    -200, 
    -215.309112548828, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -2274.43896484375, 
    -2058.82666015625, 
    -1128.07666015625, 
    -641.117614746094, 
    -145.055236816406, 
    -109.227256774902, 
    -103.238059997559, 
    -127.018707275391, 
    -237.283081054688, 
    52.9443969726562, 
    56.6110687255859, 
    496.511108398438, 
    1064.53332519531, 
    1107.31103515625, 
    1150.16943359375, 
    1003.97497558594, 
    888.469421386719, 
    874.541625976562, 
    841.388854980469, 
    879.808349609375, 
    1099.73608398438, 
    1337.375, 
    1166.322265625, 
    949.891662597656, 
    999.827758789062, 
    964.388916015625, 
    785.502746582031, 
    732.602783203125, 
    459.458343505859, 
    490.930541992188, 
    695.525024414062, 
    751.491638183594, 
    761.769470214844, 
    846.644409179688, 
    849.16943359375, 
    640.58056640625, 
    660.913879394531, 
    558.3388671875, 
    401.280548095703, 
    412.397216796875, 
    503.300018310547, 
    602.186096191406, 
    676.852783203125, 
    573.811157226562, 
    370.424987792969, 
    310.527770996094, 
    299.369445800781, 
    252.447235107422, 
    358.441680908203, 
    326.25, 
    318.113891601562, 
    330.383331298828, 
    211.29443359375, 
    83.4194488525391, 
    -81.908332824707, 
    123.570709228516, 
    272.228302001953, 
    101.846290588379, 
    31.2292079925537, 
    214.465713500977, 
    354.716186523438, 
    357.183319091797, 
    268.908355712891, 
    330.363891601562, 
    541.288879394531, 
    382.475006103516, 
    477.255554199219, 
    431.79443359375, 
    625.011108398438, 
    823.597229003906, 
    599.79443359375, 
    1077.04443359375, 
    1111.07775878906, 
    499.886108398438, 
    1448.15270996094, 
    1426.01391601562, 
    1085.54724121094, 
    956.41943359375, 
    753.702819824219, 
    460.033325195312, 
    349.616668701172, 
    356.733337402344, 
    393.558349609375, 
    427.813873291016, 
    436.561096191406, 
    348.725006103516, 
    237.447219848633, 
    254.766662597656, 
    377.427764892578, 
    382.20556640625, 
    449.422210693359, 
    487.652770996094, 
    511.45556640625, 
    456.016662597656, 
    502.983337402344, 
    381.594451904297, 
    660.677734375, 
    658.516662597656, 
    554.150024414062, 
    231.699996948242, 
    95.1472244262695, 
    202.308334350586, 
    238.541656494141, 
    83.8027801513672, 
    109.863891601562, 
    119.944442749023, 
    227.436111450195, 
    277.211120605469, 
    252.266662597656, 
    184.675003051758, 
    61.0666656494141, 
    156.552780151367, 
    169.677780151367, 
    48.277774810791, 
    64.6861114501953, 
    73.8777770996094, 
    40.3805541992188, 
    23.8999996185303, 
    -30.3444442749023, 
    312.480560302734, 
    432.713897705078, 
    437.872222900391, 
    280.783325195312, 
    239.533325195312, 
    462.555541992188, 
    1066.84997558594, 
    -23.5525760650635, 
    -391.491241455078, 
    -200, 
    -381.430816650391, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -256.145294189453, 
    -200,
  
    -2104.84545898438, 
    -1887.90502929688, 
    -383.661926269531, 
    -150.094528198242, 
    -130.391830444336, 
    -96.9208755493164, 
    -87.5234527587891, 
    -72.2585220336914, 
    -0.348558038473129, 
    136.34504699707, 
    39.5907440185547, 
    413.586120605469, 
    758.1611328125, 
    1191.177734375, 
    1180.41662597656, 
    1218.0888671875, 
    1132.39440917969, 
    1208.94445800781, 
    1137.08605957031, 
    927.136108398438, 
    920.288879394531, 
    1201.125, 
    1320.45556640625, 
    1440.95556640625, 
    1221.98059082031, 
    888.677795410156, 
    711.738891601562, 
    646.702758789062, 
    587.977783203125, 
    485.933349609375, 
    498.558349609375, 
    710.650024414062, 
    625.427795410156, 
    594.875, 
    707.799987792969, 
    718.891662597656, 
    645.536071777344, 
    649.799987792969, 
    523.027770996094, 
    437.002777099609, 
    478.027770996094, 
    506.041687011719, 
    566.852783203125, 
    439.869445800781, 
    328.183349609375, 
    232.313888549805, 
    249.241668701172, 
    324.461120605469, 
    308.441650390625, 
    211.777786254883, 
    149.355560302734, 
    156.163879394531, 
    29.3611106872559, 
    139.66389465332, 
    95.2305526733398, 
    -9.22191619873047, 
    107.985107421875, 
    113.798408508301, 
    25.2232704162598, 
    268.25830078125, 
    194.891555786133, 
    167.252777099609, 
    177.975006103516, 
    415.183349609375, 
    363.5, 
    444.161102294922, 
    503.899993896484, 
    649.924987792969, 
    468.502777099609, 
    721.155578613281, 
    619.241638183594, 
    901.647216796875, 
    309.113891601562, 
    665.597229003906, 
    1434.99169921875, 
    1274.11108398438, 
    1073.06945800781, 
    838.336120605469, 
    681.061096191406, 
    508.813873291016, 
    444.049987792969, 
    285.58056640625, 
    462.261108398438, 
    421.341674804688, 
    481.030548095703, 
    386.91943359375, 
    384.177764892578, 
    398.552764892578, 
    338.736114501953, 
    401.069427490234, 
    581.877746582031, 
    478.649993896484, 
    504.572204589844, 
    318.488891601562, 
    574.802795410156, 
    541.888916015625, 
    553.95556640625, 
    433.772216796875, 
    503.33056640625, 
    416.855560302734, 
    149.719451904297, 
    249.516662597656, 
    322.833343505859, 
    196.283340454102, 
    203.475006103516, 
    213.45832824707, 
    202.433334350586, 
    204.024993896484, 
    144.247222900391, 
    151.983337402344, 
    143.622222900391, 
    168.836120605469, 
    133.25, 
    109.919448852539, 
    99.6944427490234, 
    32.5944442749023, 
    46.2083320617676, 
    43.7666664123535, 
    317.819458007812, 
    623.272216796875, 
    567.263916015625, 
    481.411102294922, 
    325.063903808594, 
    395.627777099609, 
    760.944458007812, 
    1005.44171142578, 
    562.5263671875, 
    -429.012786865234, 
    -251.506118774414, 
    -434.940704345703, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200,
  
    -2025.66833496094, 
    -1386.14868164062, 
    -189.248504638672, 
    -136.513748168945, 
    -125.040954589844, 
    -75.0285263061523, 
    -75.1598815917969, 
    1.24696350097656, 
    141.174545288086, 
    199.645706176758, 
    332.064575195312, 
    20.1286354064941, 
    398.438873291016, 
    1272.20275878906, 
    1261.05004882812, 
    1302.75, 
    991.230529785156, 
    1049.45837402344, 
    1077.39440917969, 
    787.819458007812, 
    887.88330078125, 
    1042.11669921875, 
    1151.18884277344, 
    1090.06384277344, 
    960.79443359375, 
    677.313842773438, 
    559.858337402344, 
    621.905578613281, 
    663.736083984375, 
    575.741638183594, 
    586.486083984375, 
    610.086120605469, 
    510.825012207031, 
    456.858337402344, 
    579.783325195312, 
    644.908325195312, 
    740.172241210938, 
    748.844421386719, 
    547.027770996094, 
    487.527770996094, 
    424.030548095703, 
    383.380554199219, 
    416.672210693359, 
    288.683349609375, 
    302.097229003906, 
    256.094451904297, 
    257.350006103516, 
    291.70556640625, 
    313.594451904297, 
    215.744445800781, 
    215.20832824707, 
    7.91388893127441, 
    73.8444442749023, 
    195.905548095703, 
    163.447219848633, 
    5.47475719451904, 
    66.3642120361328, 
    142.519348144531, 
    156.29850769043, 
    247.531875610352, 
    140.1796875, 
    342.327789306641, 
    330.019439697266, 
    391.911102294922, 
    359.691680908203, 
    353.319427490234, 
    301.933319091797, 
    407.944458007812, 
    524.758361816406, 
    533.533325195312, 
    542.538879394531, 
    582.54443359375, 
    388.375, 
    843.936096191406, 
    1121.82507324219, 
    1006, 
    703.358337402344, 
    645.700012207031, 
    512.613891601562, 
    668.119445800781, 
    540.716674804688, 
    503.527770996094, 
    490.727783203125, 
    507.266662597656, 
    516.058349609375, 
    512.79443359375, 
    372.774993896484, 
    482.725006103516, 
    376.766662597656, 
    503.211120605469, 
    610.802795410156, 
    462.019439697266, 
    410.233337402344, 
    303.280548095703, 
    574.269409179688, 
    517.483337402344, 
    468.297241210938, 
    483.316680908203, 
    430.424987792969, 
    209.91667175293, 
    193.355560302734, 
    174.388885498047, 
    209.263885498047, 
    233.263885498047, 
    213.505554199219, 
    181.883331298828, 
    182.425003051758, 
    138.997222900391, 
    72.8361129760742, 
    86.908332824707, 
    81.0722198486328, 
    58.8194427490234, 
    22.0861110687256, 
    80.4861145019531, 
    33.9944458007812, 
    65.9250030517578, 
    104.549995422363, 
    246.927780151367, 
    324.866668701172, 
    380.661102294922, 
    531.708312988281, 
    329.994445800781, 
    -52.9472198486328, 
    4.1027774810791, 
    51.7222175598145, 
    121.050003051758, 
    -290.268371582031, 
    -477.375274658203, 
    -537.518249511719, 
    -545.465759277344, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -201.309753417969, 
    -205.466064453125, 
    -205.521499633789, 
    -230.09016418457,
  
    -1901.90148925781, 
    -729.761535644531, 
    -154.481506347656, 
    -123.954650878906, 
    -24.1381797790527, 
    15.622241973877, 
    469.251586914062, 
    38.0749893188477, 
    161.031326293945, 
    254.836120605469, 
    190.875793457031, 
    114.564842224121, 
    582.352783203125, 
    916.41943359375, 
    1254.75830078125, 
    1329.86938476562, 
    1016.07775878906, 
    1133.5, 
    937.788879394531, 
    562.969421386719, 
    717.563903808594, 
    1172.11108398438, 
    1001.35559082031, 
    1169.82775878906, 
    911.9638671875, 
    508.263885498047, 
    470.886108398438, 
    524.016662597656, 
    596.361083984375, 
    655.91943359375, 
    709.833312988281, 
    664.377807617188, 
    491.436126708984, 
    422.575012207031, 
    469.552764892578, 
    650.013916015625, 
    718.897216796875, 
    650.974975585938, 
    565.791687011719, 
    469.863891601562, 
    373.049987792969, 
    341.225006103516, 
    307.583343505859, 
    270.361114501953, 
    218.58610534668, 
    270.658355712891, 
    298.511108398438, 
    303.102783203125, 
    273.700012207031, 
    201.824996948242, 
    77.9222183227539, 
    80.0416641235352, 
    74.9166641235352, 
    188.433334350586, 
    133.972213745117, 
    -37.8639678955078, 
    136.210327148438, 
    -209.26611328125, 
    27.3838691711426, 
    174.006225585938, 
    286.511108398438, 
    392.54443359375, 
    476.841674804688, 
    481.219451904297, 
    520.763854980469, 
    384.338897705078, 
    422.319458007812, 
    448.222229003906, 
    461.811096191406, 
    516.844421386719, 
    596.052795410156, 
    871.408325195312, 
    731.022216796875, 
    760.319458007812, 
    959.491638183594, 
    698.783325195312, 
    681.049987792969, 
    741.5, 
    698.788879394531, 
    651.058349609375, 
    462.555541992188, 
    452.41943359375, 
    443.811126708984, 
    455.411102294922, 
    355.524993896484, 
    343.399993896484, 
    396.405548095703, 
    482.547210693359, 
    549.875, 
    671.483337402344, 
    635.369445800781, 
    485.105560302734, 
    310.008331298828, 
    349.063903808594, 
    453.922210693359, 
    398.711120605469, 
    457.680572509766, 
    567.74169921875, 
    538.41943359375, 
    236.669448852539, 
    57.6222229003906, 
    101.958335876465, 
    118.627777099609, 
    151.483337402344, 
    141.95832824707, 
    141.069442749023, 
    138.444442749023, 
    84.7777786254883, 
    80.5083312988281, 
    8.78055572509766, 
    27.1944446563721, 
    39.1333351135254, 
    40.0361099243164, 
    9.00555515289307, 
    33.5305557250977, 
    32.3722229003906, 
    90.8916625976562, 
    151.105560302734, 
    55.3583335876465, 
    262.247222900391, 
    -95.875, 
    -462.380554199219, 
    -334.33056640625, 
    311.816680908203, 
    670.977783203125, 
    494.408325195312, 
    472.188903808594, 
    -77.0451126098633, 
    -275.722808837891, 
    -671.353393554688, 
    -201.105712890625, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -226.569305419922, 
    -262.249114990234, 
    -236.336975097656, 
    -218.359329223633,
  
    -1748.34399414062, 
    -480.887725830078, 
    -161.479187011719, 
    -121.027328491211, 
    -34.3427734375, 
    155.175003051758, 
    343.600006103516, 
    324.577789306641, 
    999.033325195312, 
    885.25, 
    642.622253417969, 
    879.163879394531, 
    767.799987792969, 
    1193.96105957031, 
    1068.78332519531, 
    1240.4638671875, 
    1128.32775878906, 
    1151.27770996094, 
    1027.3583984375, 
    840.733337402344, 
    817.938903808594, 
    758.111083984375, 
    730.4111328125, 
    784.833312988281, 
    724.299987792969, 
    517.472229003906, 
    502.194427490234, 
    535.288879394531, 
    579.452758789062, 
    679.802795410156, 
    773.822204589844, 
    788.091674804688, 
    577.091674804688, 
    577.966674804688, 
    461.08056640625, 
    527.316650390625, 
    526.497253417969, 
    491.41943359375, 
    500.613891601562, 
    454.625, 
    359.013885498047, 
    354.225006103516, 
    347.636108398438, 
    236.611114501953, 
    220.938888549805, 
    222.363891601562, 
    253.811111450195, 
    248.322219848633, 
    193.858337402344, 
    179.300003051758, 
    171.633331298828, 
    129.41667175293, 
    64.2722244262695, 
    29.7055549621582, 
    69.9138870239258, 
    103.188888549805, 
    30.8249988555908, 
    -1.03333330154419, 
    49.0305557250977, 
    163.890197753906, 
    137.638885498047, 
    226.408340454102, 
    387.899993896484, 
    468.922210693359, 
    401.494445800781, 
    369.858337402344, 
    404.397216796875, 
    274.752777099609, 
    369.286102294922, 
    483.236114501953, 
    533.811096191406, 
    737.808349609375, 
    798.988891601562, 
    682.241638183594, 
    666.447204589844, 
    790.486145019531, 
    736.825012207031, 
    768.380554199219, 
    683.158325195312, 
    544.622253417969, 
    412.733337402344, 
    400.616668701172, 
    407.600006103516, 
    418.941680908203, 
    375.186126708984, 
    310.408325195312, 
    423.625, 
    464.266662597656, 
    556.897216796875, 
    632.969482421875, 
    680.458312988281, 
    416.583343505859, 
    299.116668701172, 
    342.336120605469, 
    341.452789306641, 
    334.369445800781, 
    529.844421386719, 
    605.505554199219, 
    381.450012207031, 
    176.972229003906, 
    25.8138885498047, 
    60.091667175293, 
    122.269439697266, 
    183.636108398438, 
    64.8694458007812, 
    57.663890838623, 
    76.9416656494141, 
    49.625, 
    15.8361110687256, 
    9.75833320617676, 
    -60.936107635498, 
    2.69444441795349, 
    45.4777755737305, 
    45.1222229003906, 
    42.8388900756836, 
    62.3805541992188, 
    38.0694465637207, 
    40.5027770996094, 
    -22.4388885498047, 
    -84.125, 
    -214, 
    -140.744445800781, 
    349.841674804688, 
    269.694458007812, 
    713.902770996094, 
    362.594451904297, 
    732.102783203125, 
    276.430541992188, 
    247.649993896484, 
    81.8329162597656, 
    -469.679351806641, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -250.989181518555, 
    -266.704711914062, 
    -231.11506652832, 
    -211.753372192383, 
    -207.15998840332,
  
    -1145.51843261719, 
    -840.685913085938, 
    -161.523132324219, 
    -83.1260986328125, 
    60.7058334350586, 
    797.408325195312, 
    784.577819824219, 
    752.802795410156, 
    510.702789306641, 
    1275.10827636719, 
    1060.11108398438, 
    1243.46948242188, 
    1334.27221679688, 
    1567.302734375, 
    1270.47229003906, 
    1769.09167480469, 
    1182.81945800781, 
    1271.02783203125, 
    1184.67492675781, 
    974.877807617188, 
    1125.03051757812, 
    1122.86108398438, 
    1023.11389160156, 
    974.79443359375, 
    675.772216796875, 
    466.936096191406, 
    570.736145019531, 
    640.538879394531, 
    528.452758789062, 
    630.849975585938, 
    793.691650390625, 
    731.29443359375, 
    713.54443359375, 
    664.177795410156, 
    517.872192382812, 
    436.736114501953, 
    307.83056640625, 
    364.055572509766, 
    382.983337402344, 
    375.305572509766, 
    292.808349609375, 
    229.691665649414, 
    368.858337402344, 
    233.122222900391, 
    232.705551147461, 
    192.875, 
    177.625, 
    205.713882446289, 
    60.8833312988281, 
    170.238891601562, 
    116.927780151367, 
    42.2194442749023, 
    3.77777814865112, 
    5.52222204208374, 
    43.8472213745117, 
    122.886108398438, 
    167.013885498047, 
    119.14722442627, 
    2.94444465637207, 
    -59.5111083984375, 
    -0.405555784702301, 
    190.297225952148, 
    253.438888549805, 
    309.450012207031, 
    286.141662597656, 
    320.033325195312, 
    334.994445800781, 
    260.383331298828, 
    304.125, 
    334.255554199219, 
    406.897216796875, 
    538.319458007812, 
    533.113891601562, 
    497.161102294922, 
    571.452758789062, 
    717.688903808594, 
    779.0888671875, 
    743.802795410156, 
    650.630554199219, 
    507.102783203125, 
    415.755554199219, 
    379.933319091797, 
    352.105560302734, 
    342.183349609375, 
    350.924987792969, 
    321.841674804688, 
    316.688873291016, 
    320.566680908203, 
    456.436096191406, 
    505.697235107422, 
    544.436096191406, 
    470.361114501953, 
    365.119445800781, 
    346.25, 
    498.077789306641, 
    310.238891601562, 
    353.577789306641, 
    255.227783203125, 
    149.449996948242, 
    169.319442749023, 
    88.2055511474609, 
    156.180557250977, 
    145.58610534668, 
    66.5166625976562, 
    25.6444454193115, 
    -3.45000004768372, 
    -13.3722219467163, 
    -30.286111831665, 
    -83.1305541992188, 
    -42.1166648864746, 
    -9.90277767181396, 
    13.3138885498047, 
    -43.1361122131348, 
    7.2722225189209, 
    46.7944450378418, 
    66.4305572509766, 
    35.6777763366699, 
    -6.52500009536743, 
    -84.7888870239258, 
    -153.944442749023, 
    63.1861114501953, 
    385.313903808594, 
    548.597229003906, 
    530.130554199219, 
    671.825012207031, 
    571.83056640625, 
    602.174987792969, 
    330.144439697266, 
    228.677780151367, 
    -302.822875976562, 
    -438.626098632812, 
    -213.450103759766, 
    -200, 
    -251.863098144531, 
    -200, 
    -200, 
    -200, 
    -200, 
    -246.625305175781, 
    -258.931976318359, 
    -228.884368896484,
  
    -984.08740234375, 
    -218.98860168457, 
    -158.999404907227, 
    215.511260986328, 
    443.91943359375, 
    415.43212890625, 
    1340.74719238281, 
    1207.49450683594, 
    1386.63061523438, 
    1737.33618164062, 
    1765.71948242188, 
    1802.12780761719, 
    1709.27502441406, 
    1594.01672363281, 
    1453.62219238281, 
    1625.67224121094, 
    1010.51391601562, 
    1197.39721679688, 
    1286.13610839844, 
    1078.88330078125, 
    1226.03051757812, 
    1267.91662597656, 
    1288.63891601562, 
    872.077758789062, 
    536.797241210938, 
    608.383361816406, 
    720.686096191406, 
    691.030578613281, 
    417.899993896484, 
    670.886108398438, 
    800.325012207031, 
    845.941650390625, 
    879.075012207031, 
    676.116638183594, 
    523.733337402344, 
    470.344451904297, 
    420.758331298828, 
    371.319458007812, 
    358.486114501953, 
    273.302764892578, 
    239.46110534668, 
    198.558334350586, 
    199.477783203125, 
    238.125, 
    186.655548095703, 
    149.774993896484, 
    143.969451904297, 
    121.025001525879, 
    100.683334350586, 
    113.666664123535, 
    105.35555267334, 
    43.0388870239258, 
    88.2722244262695, 
    -284.438873291016, 
    -111.419441223145, 
    157.505554199219, 
    44.0388870239258, 
    -88.1972198486328, 
    76.3388900756836, 
    51.8194427490234, 
    19.0722217559814, 
    83.2916641235352, 
    113.158332824707, 
    109.908332824707, 
    195.25, 
    228.847229003906, 
    141.497222900391, 
    12.0749998092651, 
    134.822219848633, 
    512.488891601562, 
    450.569458007812, 
    446.322235107422, 
    295.800018310547, 
    295.700012207031, 
    514.219421386719, 
    680.738891601562, 
    763.933349609375, 
    848.886108398438, 
    579.261108398438, 
    380.863891601562, 
    315.252777099609, 
    329.391662597656, 
    338.597229003906, 
    369.894439697266, 
    332.727783203125, 
    315.413879394531, 
    236.074996948242, 
    247.324996948242, 
    343.416656494141, 
    369.766662597656, 
    378.172210693359, 
    439.741668701172, 
    422.619445800781, 
    472.2861328125, 
    461.555541992188, 
    286.899993896484, 
    258.377777099609, 
    212.363891601562, 
    122.077774047852, 
    100.050003051758, 
    91.0388870239258, 
    111.908332824707, 
    127.019439697266, 
    17.2611103057861, 
    -4.21111106872559, 
    -16.1555557250977, 
    -47.3472213745117, 
    -61.5777778625488, 
    -60.4722213745117, 
    -39.591667175293, 
    -29.2722225189209, 
    -67.908332824707, 
    -120.122222900391, 
    -21.3111114501953, 
    26.6500015258789, 
    82.4055557250977, 
    103.436111450195, 
    4.37777805328369, 
    -168.877777099609, 
    -128.147216796875, 
    326.877777099609, 
    484.325012207031, 
    498.813903808594, 
    569.597229003906, 
    880.155578613281, 
    766.536071777344, 
    212.255554199219, 
    365.724090576172, 
    332.438903808594, 
    298.674987792969, 
    -426.7900390625, 
    -401.512878417969, 
    -202.291564941406, 
    -200, 
    -200, 
    -200, 
    -200, 
    -200, 
    -229.111099243164, 
    -271.193603515625, 
    -284.998687744141,
  
    -1002.51446533203, 
    -216.593414306641, 
    -143.20930480957, 
    67.745964050293, 
    408.697235107422, 
    905.016662597656, 
    876.305541992188, 
    729.694458007812, 
    1672.97778320312, 
    1750.66943359375, 
    1813.052734375, 
    1845.14721679688, 
    1714.41943359375, 
    1536.33337402344, 
    1247.18615722656, 
    1149.29443359375, 
    1031.56384277344, 
    1121.55834960938, 
    1232.33056640625, 
    1206.28894042969, 
    1389.38061523438, 
    1207.32214355469, 
    1441.13891601562, 
    1187.34729003906, 
    674.761108398438, 
    835.158325195312, 
    891.027770996094, 
    772.083312988281, 
    614.119445800781, 
    770.33056640625, 
    718.027770996094, 
    936.7861328125, 
    853.5, 
    522.722229003906, 
    619.313903808594, 
    456.322235107422, 
    305.763885498047, 
    431.941680908203, 
    444.924987792969, 
    358.541656494141, 
    215.08610534668, 
    138.677780151367, 
    133.019439697266, 
    165.044448852539, 
    142.633331298828, 
    108.955558776855, 
    120.155555725098, 
    86.6388931274414, 
    -28.8694438934326, 
    31.5944442749023, 
    63.6777801513672, 
    76.6944427490234, 
    65.4138870239258, 
    -1.65277874469757, 
    -225.755554199219, 
    37.5583343505859, 
    0.975000083446503, 
    -69.7666625976562, 
    4.89444446563721, 
    88.0166625976562, 
    4.66944456100464, 
    -93.7555541992188, 
    129.033340454102, 
    142.636108398438, 
    182.227767944336, 
    181.861114501953, 
    134.061111450195, 
    231.577774047852, 
    216.919448852539, 
    480.763885498047, 
    496.063903808594, 
    448.549987792969, 
    371.605560302734, 
    373.244445800781, 
    467.386108398438, 
    630.633361816406, 
    583.530578613281, 
    538.813903808594, 
    382.430541992188, 
    224.927780151367, 
    234.891662597656, 
    192.661117553711, 
    260.166656494141, 
    288.591674804688, 
    217.074996948242, 
    217.752777099609, 
    211.477783203125, 
    151.230545043945, 
    252.588882446289, 
    296.133331298828, 
    351.108337402344, 
    404.424987792969, 
    370.794464111328, 
    395.155548095703, 
    392.061096191406, 
    356.522216796875, 
    255.886108398438, 
    192.672225952148, 
    107.14722442627, 
    63.3583335876465, 
    11.4305553436279, 
    31.2666664123535, 
    -23.0944442749023, 
    -35.7027778625488, 
    -66.6833343505859, 
    -68.5027770996094, 
    -74.2472229003906, 
    -82.1222229003906, 
    -65.25, 
    -51.7249984741211, 
    -132.786102294922, 
    -157.080551147461, 
    -94.3472213745117, 
    -50.0416679382324, 
    4.91388893127441, 
    57.4916648864746, 
    110.783332824707, 
    110.519439697266, 
    -10.5250005722046, 
    220.050003051758, 
    202.661102294922, 
    542.936096191406, 
    395.780548095703, 
    726.708312988281, 
    901.155517578125, 
    928.436096191406, 
    626.783325195312, 
    426.308349609375, 
    496.899993896484, 
    518.474975585938, 
    -309.54248046875, 
    -440.347991943359, 
    -193.103790283203, 
    -197.212066650391, 
    -200, 
    -200, 
    -200, 
    -200, 
    -251.166259765625, 
    -384.484039306641, 
    -521.699157714844,
  
    -1078.08142089844, 
    -348.781219482422, 
    -163.176513671875, 
    -85.9037094116211, 
    501.538879394531, 
    865.738891601562, 
    530.655578613281, 
    226.078857421875, 
    767.561096191406, 
    978.611083984375, 
    799.961120605469, 
    1215.81665039062, 
    1579.18884277344, 
    1780.19995117188, 
    1466.75830078125, 
    1472.43054199219, 
    941.49169921875, 
    1128.55834960938, 
    1449.52783203125, 
    1133.15563964844, 
    1393.23889160156, 
    1576.47229003906, 
    1626.125, 
    1026.84997558594, 
    954.586120605469, 
    978.627746582031, 
    925.130554199219, 
    690.444458007812, 
    772.302795410156, 
    780.855529785156, 
    615.780517578125, 
    853.444458007812, 
    756.591674804688, 
    893.844421386719, 
    649.761108398438, 
    335.605560302734, 
    460.258331298828, 
    538.727783203125, 
    542.66943359375, 
    329.369445800781, 
    233.405563354492, 
    163.150009155273, 
    129.952774047852, 
    154.524993896484, 
    131.925003051758, 
    133.597229003906, 
    156.425003051758, 
    155.46110534668, 
    155.08610534668, 
    68.091667175293, 
    53.2305526733398, 
    62.1166648864746, 
    47.8472213745117, 
    -93.5083312988281, 
    -11.5083332061768, 
    234.591659545898, 
    -15.152777671814, 
    -93.1555557250977, 
    -191.508331298828, 
    -141.602783203125, 
    30.5, 
    -101.963882446289, 
    231, 
    226.422225952148, 
    185.213897705078, 
    193.699996948242, 
    248.5, 
    351.022216796875, 
    290.638885498047, 
    328.863891601562, 
    381.088897705078, 
    347.511108398438, 
    316.188873291016, 
    264.822235107422, 
    340.725006103516, 
    358.422210693359, 
    387.125, 
    340.336120605469, 
    308.533325195312, 
    231.400009155273, 
    255.619445800781, 
    158.991668701172, 
    165.991668701172, 
    209.352767944336, 
    200.847229003906, 
    157.149993896484, 
    154.602783203125, 
    171.16667175293, 
    315.25, 
    373.113891601562, 
    427.180572509766, 
    337.752777099609, 
    299.155548095703, 
    303.841674804688, 
    325.469451904297, 
    324.463897705078, 
    268.261108398438, 
    186.994445800781, 
    76.0138931274414, 
    40.8722229003906, 
    22.747220993042, 
    3.8611114025116, 
    -39.1027793884277, 
    -41.4444427490234, 
    -94.3388900756836, 
    -92.3027801513672, 
    -116.372222900391, 
    -61.841667175293, 
    -66.6361083984375, 
    -56.1472206115723, 
    -91.5222244262695, 
    -116.444442749023, 
    -104.675003051758, 
    -28.8611106872559, 
    58.8638877868652, 
    81.0805511474609, 
    140.388885498047, 
    170.327774047852, 
    -60.8083343505859, 
    406.66943359375, 
    238.53889465332, 
    429.333343505859, 
    567.341674804688, 
    684.4638671875, 
    619.566650390625, 
    773, 
    597.805541992188, 
    566.9638671875, 
    462.449981689453, 
    446.405548095703, 
    -383.267456054688, 
    -464.239532470703, 
    -220.894943237305, 
    -108.85319519043, 
    -189.912460327148, 
    -200, 
    -212.603881835938, 
    -261.44482421875, 
    -304.848876953125, 
    -482.689086914062, 
    -798.920227050781,
  
    -1280.14636230469, 
    -596.089660644531, 
    -172.628768920898, 
    -149.421188354492, 
    22.0238647460938, 
    153.046890258789, 
    55.544807434082, 
    478.725006103516, 
    645.224975585938, 
    327.713897705078, 
    771.686096191406, 
    891.04443359375, 
    1051.63330078125, 
    1202.87219238281, 
    1310.56945800781, 
    1849.16662597656, 
    1168.38610839844, 
    1125.73608398438, 
    1568.52783203125, 
    1129.94165039062, 
    812.888854980469, 
    1251.15551757812, 
    1460.22778320312, 
    1270.7861328125, 
    1199.85559082031, 
    1001.9111328125, 
    787.416687011719, 
    614.4638671875, 
    851.861083984375, 
    813.872253417969, 
    975.511108398438, 
    925.533325195312, 
    883.224975585938, 
    772.308349609375, 
    473.930572509766, 
    325.183319091797, 
    392.041656494141, 
    521.880554199219, 
    513.599975585938, 
    375.572235107422, 
    255.75, 
    235.658340454102, 
    134.941665649414, 
    115.180557250977, 
    170.491668701172, 
    166.005554199219, 
    166.155563354492, 
    170.761108398438, 
    125.441665649414, 
    73.3694458007812, 
    55.5722236633301, 
    41.3138885498047, 
    -8.38333320617676, 
    -75.3555603027344, 
    24.1555557250977, 
    14.0249996185303, 
    41.6749992370605, 
    -9.81111145019531, 
    -189.205551147461, 
    15.277777671814, 
    84.5055541992188, 
    31.7361106872559, 
    115.108337402344, 
    73.9555587768555, 
    -27.2722225189209, 
    -38.1277770996094, 
    173.147216796875, 
    247.077774047852, 
    251.580551147461, 
    177.791656494141, 
    317.861114501953, 
    215.119445800781, 
    265.380554199219, 
    263.858337402344, 
    254.258331298828, 
    202.675003051758, 
    270.672241210938, 
    246.061111450195, 
    302.508331298828, 
    225.411117553711, 
    226.955551147461, 
    133.722213745117, 
    91.3694458007812, 
    168.41943359375, 
    206.180557250977, 
    109.466667175293, 
    174.641662597656, 
    276.569458007812, 
    303.666687011719, 
    302.733337402344, 
    271.799987792969, 
    153.266662597656, 
    142.058334350586, 
    146.533340454102, 
    222.597229003906, 
    255.597229003906, 
    196.122222900391, 
    145.647216796875, 
    94.6138916015625, 
    35.5750007629395, 
    -40.0555534362793, 
    -50.9555549621582, 
    -88.1861114501953, 
    -115.983329772949, 
    -141.819442749023, 
    -123.180557250977, 
    -174.411102294922, 
    -124.086112976074, 
    -95, 
    -97.158332824707, 
    -85.6638870239258, 
    -89.7722244262695, 
    -30.9416675567627, 
    28.6416664123535, 
    55.2805557250977, 
    142.666656494141, 
    219.391662597656, 
    271.058349609375, 
    102.369445800781, 
    194.127777099609, 
    234.769454956055, 
    267.694458007812, 
    265.922210693359, 
    393.683319091797, 
    651.825012207031, 
    136.483337402344, 
    495.040771484375, 
    497.504180908203, 
    372.338897705078, 
    615.108337402344, 
    -163.923980712891, 
    -472.401397705078, 
    -406.435241699219, 
    -168.713256835938, 
    -147.633666992188, 
    -196.677032470703, 
    -252.917892456055, 
    -317.878265380859, 
    -448.333221435547, 
    -597.7802734375, 
    -1102.00231933594,
  
    -1455.796875, 
    -975.036804199219, 
    -257.051635742188, 
    -187.938598632812, 
    -163.31428527832, 
    -171.281753540039, 
    -144.765289306641, 
    50.4523277282715, 
    350.750518798828, 
    556.561096191406, 
    212.290008544922, 
    725.558349609375, 
    1006.29998779297, 
    579.933349609375, 
    1050.90002441406, 
    1139.447265625, 
    1334.26110839844, 
    886.683349609375, 
    1044.57775878906, 
    901.908325195312, 
    945.777770996094, 
    1390.69714355469, 
    1283.43884277344, 
    1284.81396484375, 
    1331.81665039062, 
    1272.91394042969, 
    1082.76391601562, 
    1033.34167480469, 
    1035.76110839844, 
    1003.13610839844, 
    1015.40557861328, 
    951.394470214844, 
    676.613891601562, 
    486.002777099609, 
    642.547241210938, 
    447.019439697266, 
    294.694427490234, 
    481.536102294922, 
    558.913879394531, 
    507.549987792969, 
    280.100006103516, 
    159.70832824707, 
    148.79167175293, 
    140.136108398438, 
    140.191665649414, 
    107.127777099609, 
    168.155548095703, 
    183.372222900391, 
    90.7555541992188, 
    -16.8611106872559, 
    10.5361108779907, 
    34.7027778625488, 
    86.8583297729492, 
    -38.494441986084, 
    -27.6638889312744, 
    -57.2416687011719, 
    -9.00555515289307, 
    -57.6944427490234, 
    -139.899993896484, 
    38.2277755737305, 
    -92.125, 
    -47.4305534362793, 
    41.8055572509766, 
    -48.7277793884277, 
    -164.155548095703, 
    -168.622222900391, 
    24.9972229003906, 
    108.805557250977, 
    177.355545043945, 
    268.497222900391, 
    296.5888671875, 
    239.138885498047, 
    180.725006103516, 
    143.169448852539, 
    152.494445800781, 
    172.511108398438, 
    182.449996948242, 
    169.547225952148, 
    167.830551147461, 
    178.158340454102, 
    208.016662597656, 
    107.358337402344, 
    90.0277786254883, 
    107.016662597656, 
    115.830551147461, 
    58.5555572509766, 
    218.947219848633, 
    297.350006103516, 
    263.674987792969, 
    175.722229003906, 
    111.236114501953, 
    166.927780151367, 
    94.2777786254883, 
    9.86388874053955, 
    217.636108398438, 
    176.941665649414, 
    50.9305572509766, 
    158.033325195312, 
    53.3138885498047, 
    -31.6361103057861, 
    -71.966667175293, 
    -89.2583312988281, 
    -194.505554199219, 
    -115.572219848633, 
    -140.330551147461, 
    -176.747222900391, 
    -172.786117553711, 
    -179.619445800781, 
    -127.791664123535, 
    -79.875, 
    -47.6777763366699, 
    -24.3555564880371, 
    -4.38888883590698, 
    101.913887023926, 
    138.422225952148, 
    217.66389465332, 
    330.975006103516, 
    237.666656494141, 
    45.9583320617676, 
    362.386108398438, 
    399.588897705078, 
    589.016662597656, 
    599.469421386719, 
    678.380554199219, 
    775.744445800781, 
    1034.85559082031, 
    814.152770996094, 
    303.355560302734, 
    71.9504623413086, 
    500.679809570312, 
    -255.793487548828, 
    -493.922210693359, 
    -495.302551269531, 
    -278.800598144531, 
    -224.276214599609, 
    -235.938568115234, 
    -276.640899658203, 
    -316.463989257812, 
    -390.670166015625, 
    -552.245178222656, 
    -1100.72998046875,
  
    -1904.20629882812, 
    -1635.94348144531, 
    -609.961853027344, 
    -213.003204345703, 
    -185.80696105957, 
    -206.049453735352, 
    -269.835327148438, 
    -189.124481201172, 
    -189.766403198242, 
    -103.195365905762, 
    -68.6347427368164, 
    31.0535488128662, 
    376.08056640625, 
    659.086120605469, 
    464.602752685547, 
    810.519470214844, 
    904.522216796875, 
    884.552795410156, 
    200.622222900391, 
    233.05322265625, 
    897.905578613281, 
    1048.39440917969, 
    1674.17504882812, 
    1625.30834960938, 
    1340.80554199219, 
    1588.58056640625, 
    1218.52502441406, 
    1179.54162597656, 
    1370.39172363281, 
    1321.06945800781, 
    927.099975585938, 
    1112.06665039062, 
    851.611083984375, 
    755.430541992188, 
    814.711120605469, 
    519.913879394531, 
    403.197235107422, 
    544.833312988281, 
    682.125, 
    364.991668701172, 
    213.183334350586, 
    144.469436645508, 
    108.47777557373, 
    134.938888549805, 
    172.480560302734, 
    193.305557250977, 
    179.658340454102, 
    188.25, 
    101.261108398438, 
    72.5305557250977, 
    25.1527767181396, 
    -34.1861114501953, 
    -146.783340454102, 
    -59.8833351135254, 
    -151.350006103516, 
    -101.441665649414, 
    -73.1611099243164, 
    -163.730560302734, 
    -135.294448852539, 
    31.3527774810791, 
    -63.7777786254883, 
    -103.047218322754, 
    96.7138900756836, 
    43.125, 
    -73.6388854980469, 
    -51.9777755737305, 
    15.2194442749023, 
    56.6027793884277, 
    117.088890075684, 
    169.855560302734, 
    236.024993896484, 
    226.002777099609, 
    99.6222229003906, 
    32.8472213745117, 
    72.0388870239258, 
    125.213890075684, 
    98.1305541992188, 
    62.4361114501953, 
    79.3499984741211, 
    127.386108398438, 
    76.9416656494141, 
    55.9611129760742, 
    60.7583351135254, 
    46.8638877868652, 
    94.5555572509766, 
    51.283332824707, 
    83.1833343505859, 
    176.730560302734, 
    167.780548095703, 
    137.161117553711, 
    185.08332824707, 
    161.472229003906, 
    117.194442749023, 
    91.033332824707, 
    150.527770996094, 
    56.3722229003906, 
    -103.677772521973, 
    133.941665649414, 
    30.9611110687256, 
    -95.6027755737305, 
    13.1611108779907, 
    -93.9499969482422, 
    -127.847221374512, 
    -140.094451904297, 
    -148.627777099609, 
    -115.094444274902, 
    -154.775009155273, 
    -198.861114501953, 
    -233.074996948242, 
    -80.2444458007812, 
    9.26388931274414, 
    -21.0611114501953, 
    23.4277782440186, 
    -45.2388877868652, 
    -135.561111450195, 
    -72.6722259521484, 
    34.6333312988281, 
    7.79722261428833, 
    262.45556640625, 
    431.963897705078, 
    499.658325195312, 
    500.961120605469, 
    531.724975585938, 
    627.402770996094, 
    675.850036621094, 
    576.594421386719, 
    279.113891601562, 
    -13.0972118377686, 
    -89.3597869873047, 
    -213.382202148438, 
    -521.917663574219, 
    -686.404602050781, 
    -476.9560546875, 
    -410.858154296875, 
    -305.535034179688, 
    -281.026947021484, 
    -289.068817138672, 
    -303.296478271484, 
    -313.916229248047, 
    -378.286468505859, 
    -1071.47680664062,
  
    -1995.84436035156, 
    -1816.19177246094, 
    -1724.7578125, 
    -1362.40075683594, 
    -475.337768554688, 
    -344.816070556641, 
    -196.469253540039, 
    -232.626525878906, 
    -404.350677490234, 
    -245.577484130859, 
    -273.357879638672, 
    -195.303756713867, 
    -199.969390869141, 
    113.609077453613, 
    361.297882080078, 
    396.327789306641, 
    391.691925048828, 
    262.823974609375, 
    473.44970703125, 
    16.4071559906006, 
    320.575012207031, 
    1106.21118164062, 
    1307.57495117188, 
    898.083312988281, 
    1590.60559082031, 
    1641.95007324219, 
    1392.73059082031, 
    1101.93615722656, 
    1390.04174804688, 
    1216.177734375, 
    943.400024414062, 
    1013.37780761719, 
    970.130554199219, 
    929.658325195312, 
    518.752807617188, 
    536.958312988281, 
    593.488891601562, 
    568.66943359375, 
    523.541687011719, 
    453.502777099609, 
    334.75, 
    162.886108398438, 
    107.172225952148, 
    312.680541992188, 
    197.21110534668, 
    93.5944442749023, 
    149.430557250977, 
    132.088882446289, 
    144.272216796875, 
    164.175003051758, 
    59.6944427490234, 
    -42.0666656494141, 
    -133.091674804688, 
    -145.822219848633, 
    -58.0805549621582, 
    -14.222222328186, 
    -40.4000015258789, 
    -133.722229003906, 
    -90.7750015258789, 
    -50.2805557250977, 
    -46.341667175293, 
    -18.75, 
    23.8166656494141, 
    68.5527801513672, 
    24.0694446563721, 
    16.7583332061768, 
    27.4027786254883, 
    2.7138888835907, 
    75.783332824707, 
    132.274993896484, 
    109.783332824707, 
    83.7305526733398, 
    16.7055549621582, 
    -42.6166648864746, 
    -13.8805551528931, 
    68.8222198486328, 
    61.586109161377, 
    -69.3555526733398, 
    -33.8166656494141, 
    14.7555561065674, 
    -13.8333330154419, 
    23.4555549621582, 
    22.8166656494141, 
    42.9777793884277, 
    48.9777755737305, 
    38.6333312988281, 
    32.8805541992188, 
    76.4861145019531, 
    115.347221374512, 
    134.53889465332, 
    124.005554199219, 
    80.1944427490234, 
    62.9638900756836, 
    28.3083343505859, 
    -2.98055553436279, 
    -36.1388893127441, 
    -20.6388893127441, 
    -41.0277786254883, 
    -9.41388893127441, 
    -67.1388854980469, 
    -45.5805549621582, 
    -172.938888549805, 
    -97.4444427490234, 
    -164.741668701172, 
    -169.224990844727, 
    -90.1222229003906, 
    -145.986114501953, 
    -123.188888549805, 
    -138.21110534668, 
    -87.9277725219727, 
    -41.0388870239258, 
    -24.033332824707, 
    -10.0138883590698, 
    15.1944437026978, 
    112.641670227051, 
    257.055572509766, 
    126.261108398438, 
    221.591674804688, 
    182.586120605469, 
    320.202758789062, 
    496.833343505859, 
    399.861114501953, 
    64.2361145019531, 
    -248.758346557617, 
    -250.680541992188, 
    -226.486114501953, 
    -42.8722267150879, 
    262.700775146484, 
    383.866668701172, 
    647.906799316406, 
    21.9704895019531, 
    -692.797119140625, 
    -494.28564453125, 
    -400.376647949219, 
    -363.573181152344, 
    -303.014556884766, 
    -294.700164794922, 
    -289.213684082031, 
    -326.503997802734, 
    -487.456787109375, 
    -994.150634765625,
  
    -2192.43627929688, 
    -2008.31298828125, 
    -1873.09924316406, 
    -1780.07080078125, 
    -1668.7041015625, 
    -1459.11450195312, 
    -1191.11730957031, 
    -826.282958984375, 
    -280.918334960938, 
    -207.792846679688, 
    -439.796905517578, 
    -366.471923828125, 
    -213.07453918457, 
    -185.271560668945, 
    -74.6026382446289, 
    -140.157409667969, 
    -96.6534423828125, 
    -99.447868347168, 
    -91.7905120849609, 
    19.8779182434082, 
    579.708312988281, 
    293.673400878906, 
    385.875, 
    1114.36669921875, 
    1177.822265625, 
    1380.88061523438, 
    1301.23889160156, 
    912.38330078125, 
    985.305541992188, 
    886.058349609375, 
    1006.69171142578, 
    672.605529785156, 
    920.33056640625, 
    949.638916015625, 
    329.891662597656, 
    559.405578613281, 
    450.683319091797, 
    451.04443359375, 
    337.947235107422, 
    259.980560302734, 
    263.011108398438, 
    217.130554199219, 
    227.683334350586, 
    396.630554199219, 
    282.394439697266, 
    257.822235107422, 
    176.074996948242, 
    95.1388931274414, 
    175.28889465332, 
    134.686111450195, 
    33.2611122131348, 
    -8.38611125946045, 
    -98.2666625976562, 
    -183.397216796875, 
    -70.8361129760742, 
    -72.5083312988281, 
    -82.0749969482422, 
    -59.8888893127441, 
    -13.7555551528931, 
    17.0222225189209, 
    32.7222213745117, 
    12.4583330154419, 
    51.3972244262695, 
    54.3333320617676, 
    9.59444427490234, 
    20.4972229003906, 
    18.4694442749023, 
    44.6722221374512, 
    99.1750030517578, 
    103.122222900391, 
    70.2583312988281, 
    35.0138893127441, 
    -38.2305564880371, 
    -93.0805511474609, 
    -64.1138916015625, 
    -17.6944446563721, 
    -42.5638885498047, 
    -118.052780151367, 
    -142.061111450195, 
    -120.908332824707, 
    -104.872222900391, 
    -117.700004577637, 
    -67.4250030517578, 
    -57.4500007629395, 
    -23.5638885498047, 
    6.6027774810791, 
    20.1416664123535, 
    57.7722206115723, 
    62.9916687011719, 
    81.3194427490234, 
    70.7583312988281, 
    -39.1388893127441, 
    -78.8000030517578, 
    -112.655555725098, 
    -118.649993896484, 
    -108.199996948242, 
    -137.608337402344, 
    -67.8333358764648, 
    -64.4055557250977, 
    -124.130554199219, 
    -217.655563354492, 
    -44.0555572509766, 
    -70.0999984741211, 
    -142.630554199219, 
    -157.730560302734, 
    -152.633331298828, 
    -154.669448852539, 
    -102.183334350586, 
    -120.47777557373, 
    -143.019439697266, 
    -127.138893127441, 
    -66.6472244262695, 
    -80.3722229003906, 
    56.5805587768555, 
    123.430557250977, 
    147.680557250977, 
    123.030555725098, 
    175.074996948242, 
    167.427780151367, 
    217.627777099609, 
    447.411102294922, 
    408.363891601562, 
    144.202774047852, 
    475.697204589844, 
    613.344421386719, 
    616.25830078125, 
    532.369445800781, 
    502.997222900391, 
    293.305572509766, 
    658.510070800781, 
    -351.056732177734, 
    -130.314010620117, 
    -399.970825195312, 
    -430.430450439453, 
    -415.124969482422, 
    -346.815399169922, 
    -302.476501464844, 
    -293.273986816406, 
    -309.353820800781, 
    -389.919097900391, 
    -802.815979003906,
  
    -2314.22875976562, 
    -2186.69555664062, 
    -2013.81372070312, 
    -1886.59997558594, 
    -2003.89123535156, 
    -1814.5576171875, 
    -1683.37231445312, 
    -1735.21875, 
    -1606.61889648438, 
    -1293.09216308594, 
    -730.59326171875, 
    -222.01579284668, 
    -203.342071533203, 
    -257.40478515625, 
    -261.014770507812, 
    -218.241928100586, 
    -402.812866210938, 
    -264.011566162109, 
    -539.002197265625, 
    -122.857284545898, 
    130.28254699707, 
    213.238891601562, 
    718.483337402344, 
    450.505554199219, 
    369.266662597656, 
    978.822204589844, 
    736.727783203125, 
    1051.697265625, 
    687.497192382812, 
    910.4638671875, 
    985.20556640625, 
    978.772216796875, 
    1256.61669921875, 
    506.602783203125, 
    538.66943359375, 
    450.013885498047, 
    423.211120605469, 
    401.005554199219, 
    344.058349609375, 
    368.20556640625, 
    339.424987792969, 
    167.058334350586, 
    140.649993896484, 
    192.197219848633, 
    192.397216796875, 
    168.997222900391, 
    125.916664123535, 
    204.894439697266, 
    55.2277793884277, 
    148.016662597656, 
    94.7611083984375, 
    70.875, 
    36.4249992370605, 
    -135.649993896484, 
    -95.7138900756836, 
    -174.96110534668, 
    -156.844451904297, 
    -64.0722198486328, 
    -9.6694450378418, 
    45.1638870239258, 
    74.9222183227539, 
    79.4166717529297, 
    76.569450378418, 
    27.9249992370605, 
    1.13333332538605, 
    37.5194435119629, 
    -39.6222229003906, 
    -22.1333332061768, 
    40.375, 
    95.2472229003906, 
    49.8972206115723, 
    8.86388874053955, 
    -42.5, 
    -55.7555541992188, 
    -68.7944412231445, 
    -149.866668701172, 
    72.7388916015625, 
    -24.0666656494141, 
    -73.7861099243164, 
    -108.097221374512, 
    -202.980560302734, 
    -311.04443359375, 
    -254.113891601562, 
    -162.233337402344, 
    -50.3972244262695, 
    -25.5194435119629, 
    -21.9972229003906, 
    3.14444446563721, 
    -9.43055534362793, 
    -26.7000007629395, 
    -82.875, 
    -117.802780151367, 
    -103.533332824707, 
    -93.9749984741211, 
    -97.3472213745117, 
    -137.358337402344, 
    -208.088897705078, 
    -139.761108398438, 
    -199.802780151367, 
    -55.7805557250977, 
    -48.6055564880371, 
    -73.3944473266602, 
    -101.741668701172, 
    -120.402778625488, 
    -290.611114501953, 
    -144.138885498047, 
    -105.336112976074, 
    -79.591667175293, 
    -112.516662597656, 
    -167.050003051758, 
    -143.508331298828, 
    -80.5888900756836, 
    -31.5666675567627, 
    42.0611114501953, 
    121.974998474121, 
    97.0583343505859, 
    91.283332824707, 
    137.336120605469, 
    318.866668701172, 
    477.786102294922, 
    400.861114501953, 
    408.972229003906, 
    549.983337402344, 
    433.333343505859, 
    469.927764892578, 
    662.424987792969, 
    279.683319091797, 
    253.149993896484, 
    -38.2358818054199, 
    -21.8137893676758, 
    -189.035003662109, 
    -23.4039535522461, 
    -162.303359985352, 
    -348.680908203125, 
    -378.665771484375, 
    -328.644439697266, 
    -299.362487792969, 
    -275.340911865234, 
    -300.470916748047, 
    -471.573608398438, 
    -1436.93078613281,
  
    -2534.9560546875, 
    -2384.49877929688, 
    -2220.9482421875, 
    -2175.37036132812, 
    -2058.61401367188, 
    -1882.17858886719, 
    -1826.4990234375, 
    -2020.56164550781, 
    -1921.0419921875, 
    -1713.33520507812, 
    -1720.47399902344, 
    -1332.21496582031, 
    -849.78125, 
    -314.466278076172, 
    -307.630126953125, 
    -227.866455078125, 
    -452.039093017578, 
    -474.006195068359, 
    -427.905059814453, 
    -271.404571533203, 
    -256.583312988281, 
    -98.3254699707031, 
    102.73055267334, 
    136.95832824707, 
    688.316650390625, 
    274.615966796875, 
    574.597229003906, 
    867.302795410156, 
    74.6964111328125, 
    1102.56665039062, 
    1208.05004882812, 
    990.238891601562, 
    604.216674804688, 
    563.45556640625, 
    616.722229003906, 
    399.049987792969, 
    352.288879394531, 
    299.791656494141, 
    321.286102294922, 
    181.427780151367, 
    177.233337402344, 
    215.508331298828, 
    275.413879394531, 
    235.194442749023, 
    197.844436645508, 
    134.063888549805, 
    58.1611099243164, 
    78.0722198486328, 
    -12.1694440841675, 
    -7.90000009536743, 
    -5.24722194671631, 
    40.0750007629395, 
    187.027770996094, 
    -61.8694458007812, 
    5.34166717529297, 
    -21.7277774810791, 
    -112.961112976074, 
    -71.2222213745117, 
    -24.3666667938232, 
    62.341667175293, 
    62.9416656494141, 
    -14.216667175293, 
    -1.63888907432556, 
    65.3166656494141, 
    -52.4472236633301, 
    -49.6305541992188, 
    -108.411109924316, 
    -4.65277767181396, 
    57.6305541992188, 
    46.8805541992188, 
    76.0305557250977, 
    -15.5166664123535, 
    -53.7972221374512, 
    -77.3305511474609, 
    -103.338890075684, 
    -22.6694450378418, 
    -53.5250015258789, 
    -61.1388893127441, 
    -89.8638916015625, 
    -27.2250003814697, 
    -50.5638885498047, 
    -81.7777786254883, 
    -103.741668701172, 
    -142.816665649414, 
    -55.4694442749023, 
    -78.8805541992188, 
    -108.369445800781, 
    -124.588890075684, 
    -196.230560302734, 
    -209.188888549805, 
    -111.622222900391, 
    -115.777778625488, 
    -136.027770996094, 
    -148.422210693359, 
    -183.222213745117, 
    -157.21110534668, 
    -122.880554199219, 
    -137.661102294922, 
    -160.422225952148, 
    -158.747222900391, 
    -168.525009155273, 
    -120.280555725098, 
    -156.183334350586, 
    -154.819442749023, 
    -213.355560302734, 
    -115.01944732666, 
    -52.9944458007812, 
    -49.4166641235352, 
    -73.3805541992188, 
    -88.7916641235352, 
    -89.6277770996094, 
    -95.8361129760742, 
    -30.1166667938232, 
    56.3166656494141, 
    142.786102294922, 
    192.425003051758, 
    207.936111450195, 
    189.552780151367, 
    317.163879394531, 
    426.252777099609, 
    425.763885498047, 
    572.355529785156, 
    662.211120605469, 
    677.733337402344, 
    596.997253417969, 
    562.383361816406, 
    54.564640045166, 
    -235.386611938477, 
    343.967163085938, 
    621.011108398438, 
    227.19401550293, 
    -49.0994186401367, 
    -83.6961822509766, 
    -246.115158081055, 
    -301.020416259766, 
    -275.060363769531, 
    -262.698577880859, 
    -294.321807861328, 
    -311.046417236328, 
    -1070.18579101562, 
    -2039.57775878906,
  
    -2659.52490234375, 
    -2486.11767578125, 
    -2412.181640625, 
    -2417.61059570312, 
    -2237.93725585938, 
    -2015.50720214844, 
    -2023.23266601562, 
    -2173.45727539062, 
    -1959.09521484375, 
    -2010.13110351562, 
    -1963.67944335938, 
    -1848.91979980469, 
    -1764.19750976562, 
    -1457.6611328125, 
    -1259.9912109375, 
    -520.078369140625, 
    -405.52978515625, 
    -596.726623535156, 
    -222.067016601562, 
    -203.203460693359, 
    -402.154968261719, 
    -366.819030761719, 
    -133.9150390625, 
    12.9828882217407, 
    412.549987792969, 
    720.413879394531, 
    940.055541992188, 
    230.566665649414, 
    156.768188476562, 
    1004.00280761719, 
    1090.15283203125, 
    646.602783203125, 
    259.477600097656, 
    376.149993896484, 
    593.902770996094, 
    323.263885498047, 
    348.136108398438, 
    308.930541992188, 
    224.541656494141, 
    172.302780151367, 
    271.202789306641, 
    346.799987792969, 
    334.833343505859, 
    222.613891601562, 
    221.522216796875, 
    115.094444274902, 
    147.597229003906, 
    199.661102294922, 
    105.566665649414, 
    40.9583320617676, 
    57.5472221374512, 
    13.277777671814, 
    -54.9277801513672, 
    -79.3972244262695, 
    114.76944732666, 
    -5.42500019073486, 
    -194.866668701172, 
    -55.7777786254883, 
    15.5611114501953, 
    136.636108398438, 
    26.4944458007812, 
    -88.1777801513672, 
    -0.997222125530243, 
    70.1555557250977, 
    -67.8083343505859, 
    -124.64722442627, 
    -79.2361145019531, 
    14.1388893127441, 
    50.972225189209, 
    8.63333320617676, 
    29.9527778625488, 
    -42.1722221374512, 
    -95.8250045776367, 
    -112.086112976074, 
    -86.7555541992188, 
    10.2055559158325, 
    -92.8527755737305, 
    -77.6805572509766, 
    -13.652777671814, 
    -10.4555559158325, 
    -26.4500007629395, 
    -31.2000007629395, 
    -86.3000030517578, 
    -119.258331298828, 
    -126.930557250977, 
    -153.052780151367, 
    -128.91389465332, 
    -133.936111450195, 
    -119.583335876465, 
    -123.966667175293, 
    -108.791664123535, 
    -138.277770996094, 
    -159.502777099609, 
    -157.422225952148, 
    -182.449996948242, 
    -158.688888549805, 
    -157.883331298828, 
    -180.269439697266, 
    -211.255554199219, 
    -212.475006103516, 
    -199.622222900391, 
    -176.455551147461, 
    -166.008331298828, 
    -151.71110534668, 
    -164.336120605469, 
    -84.2027816772461, 
    -97.6027755737305, 
    -94.6027755737305, 
    -110.163887023926, 
    -121.677780151367, 
    -108.308334350586, 
    -78.7944488525391, 
    -41.3444442749023, 
    17.2861099243164, 
    182.561111450195, 
    200.663879394531, 
    124.961112976074, 
    177.477783203125, 
    200.766662597656, 
    327.024993896484, 
    492.702758789062, 
    500.802764892578, 
    439.519439697266, 
    515.291687011719, 
    137.308334350586, 
    -29.4992332458496, 
    205.829177856445, 
    223.672225952148, 
    322.066650390625, 
    453.850006103516, 
    26.5268516540527, 
    16.9163112640381, 
    219.900390625, 
    -166.264785766602, 
    -261.029571533203, 
    -305.639587402344, 
    -263.772247314453, 
    -299.304962158203, 
    -353.366149902344, 
    -1310.51635742188, 
    -2211.8525390625,
  
    -2667.10766601562, 
    -2679.13623046875, 
    -2564.71313476562, 
    -2655.27856445312, 
    -2509.35180664062, 
    -2141.45654296875, 
    -2364.91723632812, 
    -2329.943359375, 
    -2134.11572265625, 
    -2220.87377929688, 
    -1894.07482910156, 
    -1905.12390136719, 
    -1836.60559082031, 
    -1779.96472167969, 
    -1777.77429199219, 
    -1593.74462890625, 
    -764.259460449219, 
    -421.54931640625, 
    -698.673034667969, 
    -1130.88037109375, 
    -494.019683837891, 
    -262.471710205078, 
    -286.168579101562, 
    -208.198760986328, 
    -66.2493515014648, 
    151.439300537109, 
    3.51937866210938, 
    244.399353027344, 
    26.3814392089844, 
    338.372772216797, 
    673.372253417969, 
    287.913879394531, 
    -35.8306427001953, 
    210.344436645508, 
    675.930541992188, 
    546.658325195312, 
    447.791656494141, 
    384.030548095703, 
    236.733337402344, 
    288.227783203125, 
    347.799987792969, 
    261.158325195312, 
    229.716659545898, 
    194.316665649414, 
    106.330551147461, 
    88.2416687011719, 
    201.530548095703, 
    280.416656494141, 
    205.147216796875, 
    39.3027763366699, 
    47.9805564880371, 
    -54.75, 
    -100.883331298828, 
    -5.22222232818604, 
    119.516670227051, 
    13.9055557250977, 
    -115.208335876465, 
    -50.6111106872559, 
    41.8444442749023, 
    66.5749969482422, 
    43.2111129760742, 
    -24.6444435119629, 
    9.09166717529297, 
    71.3944473266602, 
    74.1194458007812, 
    21.661111831665, 
    -72.2638854980469, 
    -9.11944484710693, 
    43.9000015258789, 
    31.0361099243164, 
    -37.1611099243164, 
    -72.7194442749023, 
    -112.891670227051, 
    -97.1638870239258, 
    -60.2027778625488, 
    -11.0583333969116, 
    47.6944427490234, 
    59.3722229003906, 
    39.8527793884277, 
    5.47777795791626, 
    -20.6027774810791, 
    -68.125, 
    -134.725006103516, 
    -168.29167175293, 
    -161.480560302734, 
    -174.46110534668, 
    -134.888885498047, 
    -116.366668701172, 
    -125.591667175293, 
    -137.183334350586, 
    -129.161117553711, 
    -134.95832824707, 
    -152.349990844727, 
    -114.336112976074, 
    -162.355560302734, 
    -162.752777099609, 
    -170.144439697266, 
    -197.436111450195, 
    -221.077774047852, 
    -233.902786254883, 
    -231.377777099609, 
    -203.613891601562, 
    -164.172225952148, 
    -170.436111450195, 
    -232.16667175293, 
    -109.827774047852, 
    -117.099998474121, 
    -106.60555267334, 
    -121.097221374512, 
    -163.555557250977, 
    -93.5277786254883, 
    -66.841667175293, 
    -53.6416664123535, 
    -31.9194450378418, 
    61.4000015258789, 
    111.22777557373, 
    142.5, 
    242.71110534668, 
    227.411102294922, 
    385.561126708984, 
    471.024993896484, 
    438.225006103516, 
    541.236145019531, 
    513.986083984375, 
    651.238891601562, 
    581.075012207031, 
    612.111145019531, 
    744.844421386719, 
    174.840789794922, 
    712.677795410156, 
    828.711120605469, 
    218.74560546875, 
    595.91943359375, 
    -73.7003479003906, 
    -224.685577392578, 
    -282.066131591797, 
    -277.242340087891, 
    -299.9794921875, 
    -369.966979980469, 
    -1402.17224121094, 
    -2109.42846679688,
  
    -2823.7822265625, 
    -2777.02856445312, 
    -2652.9443359375, 
    -2528.45434570312, 
    -2468.69458007812, 
    -2319.78491210938, 
    -2526.62353515625, 
    -2379.50390625, 
    -2255.7431640625, 
    -2278.34497070312, 
    -2103.28784179688, 
    -2090.45263671875, 
    -2098.4833984375, 
    -1981.82299804688, 
    -1425.22009277344, 
    -1251.203125, 
    -1404.71813964844, 
    -1643.22778320312, 
    -1642.44079589844, 
    -1556.3544921875, 
    -1596.8603515625, 
    -991.018859863281, 
    -253.032272338867, 
    -287.281463623047, 
    -326.897155761719, 
    -671.670837402344, 
    -736.778930664062, 
    -553.723693847656, 
    -77.052001953125, 
    143.65412902832, 
    -25.5112724304199, 
    -19.0725574493408, 
    96.2158126831055, 
    564.775024414062, 
    862.805541992188, 
    653.844482421875, 
    426.108337402344, 
    509.566650390625, 
    490.230560302734, 
    426.036102294922, 
    199.691665649414, 
    185.363891601562, 
    157.091659545898, 
    92.8944473266602, 
    156.969436645508, 
    139.199996948242, 
    270.244445800781, 
    412.288879394531, 
    254.813888549805, 
    60.4722213745117, 
    -12.0666675567627, 
    -28.8944435119629, 
    -75.7444458007812, 
    -0.744444370269775, 
    41.8083343505859, 
    65.9722213745117, 
    114.030555725098, 
    51.6972236633301, 
    -17.6749992370605, 
    -152.786117553711, 
    -34.533332824707, 
    -85.4555511474609, 
    -55.4555549621582, 
    54.0583343505859, 
    103.64444732666, 
    -6.47499990463257, 
    -68.1083374023438, 
    48.1138916015625, 
    15.591667175293, 
    -9.80833339691162, 
    -24.2083339691162, 
    -54.0250015258789, 
    -97.2583312988281, 
    -52.0722236633301, 
    -5.76388883590698, 
    142.419448852539, 
    103.819442749023, 
    132.449996948242, 
    105.177772521973, 
    -48.5055541992188, 
    50.4444427490234, 
    -90.0583343505859, 
    -138.705551147461, 
    -168.858337402344, 
    -180.169448852539, 
    -171.127777099609, 
    -140.486114501953, 
    -90.2611083984375, 
    -52.2583351135254, 
    -109.266670227051, 
    -116.300003051758, 
    -144.838882446289, 
    -147.994445800781, 
    -111.777778625488, 
    -165.983337402344, 
    -194.08610534668, 
    -187.619445800781, 
    -200.675003051758, 
    -231.675003051758, 
    -218.044448852539, 
    -200.547225952148, 
    -209.102783203125, 
    -165.350006103516, 
    -153.677780151367, 
    -192.763885498047, 
    -146.925003051758, 
    -124.791664123535, 
    -45.7666664123535, 
    -21.6666660308838, 
    -6.03888893127441, 
    -51.1027793884277, 
    -56.0972213745117, 
    -20.6499996185303, 
    -35.9361114501953, 
    -35.2222213745117, 
    14.402777671814, 
    67.4277801513672, 
    127.35277557373, 
    290.391662597656, 
    399.288879394531, 
    580.702758789062, 
    631.447204589844, 
    659.486145019531, 
    927.391662597656, 
    1029.81665039062, 
    915.394409179688, 
    339.836120605469, 
    348.847229003906, 
    920.472229003906, 
    1028.24169921875, 
    750.688903808594, 
    206.676513671875, 
    495.905548095703, 
    241.861114501953, 
    -152.945663452148, 
    -263.00634765625, 
    -274.658386230469, 
    -316.136413574219, 
    -436.691436767578, 
    -1443.38562011719, 
    -2070.36767578125,
  
    -2967.48608398438, 
    -2897.59130859375, 
    -2707.41796875, 
    -2615.79174804688, 
    -2516.2431640625, 
    -2507.48046875, 
    -2637.89575195312, 
    -2500.8505859375, 
    -2377.33544921875, 
    -2468.81884765625, 
    -2336.86938476562, 
    -2309.037109375, 
    -2253.5224609375, 
    -1996.7431640625, 
    -1596.89953613281, 
    -1472.25390625, 
    -1769.57360839844, 
    -1785.7939453125, 
    -1506.72705078125, 
    -1897.6259765625, 
    -1683.744140625, 
    -1551.69592285156, 
    -880.617736816406, 
    -441.976867675781, 
    -554.801696777344, 
    -276.219665527344, 
    -214.779006958008, 
    -281.850311279297, 
    -224.057144165039, 
    -201.982849121094, 
    -210.128219604492, 
    -92.2884063720703, 
    -4.92928791046143, 
    89.0103759765625, 
    387.574554443359, 
    63.2221641540527, 
    351.805541992188, 
    540.341674804688, 
    498.013885498047, 
    465.58056640625, 
    525.536071777344, 
    367.952789306641, 
    238.988891601562, 
    214.186111450195, 
    388.408325195312, 
    273.230560302734, 
    234.188888549805, 
    167.563888549805, 
    156.28889465332, 
    69.3694458007812, 
    -80.8666687011719, 
    -73.1944427490234, 
    -54.9055557250977, 
    19.6750011444092, 
    104.052780151367, 
    107.958335876465, 
    3.0722222328186, 
    44.5666656494141, 
    39.913890838623, 
    -139.066665649414, 
    -50.8666648864746, 
    -18.0499992370605, 
    -34.3388900756836, 
    -21.2638893127441, 
    -70.4694442749023, 
    -58.7583312988281, 
    -4.8972225189209, 
    162.669448852539, 
    44.0694427490234, 
    -2.3527774810791, 
    -17.4138889312744, 
    -53.158332824707, 
    -50.283332824707, 
    -31.9222221374512, 
    16.9750003814697, 
    93.6750030517578, 
    101.719444274902, 
    176.094436645508, 
    168.294448852539, 
    44.4166679382324, 
    26.7555561065674, 
    -39.2694435119629, 
    -156.397232055664, 
    -174.252777099609, 
    -168.502777099609, 
    -139.797225952148, 
    -86.3333358764648, 
    -82.0083389282227, 
    -50.9527778625488, 
    -101.927780151367, 
    -95.5777740478516, 
    -142.324996948242, 
    -118.888885498047, 
    -102.927780151367, 
    -131.133331298828, 
    -140.75, 
    -163.813888549805, 
    -134.783325195312, 
    -187.544448852539, 
    -183.491668701172, 
    -186.977767944336, 
    -198.158340454102, 
    -144.994445800781, 
    -159.011108398438, 
    -268.777770996094, 
    -239.680557250977, 
    -165.919448852539, 
    -11.1777772903442, 
    -138.441665649414, 
    -6.65833330154419, 
    -51.0222244262695, 
    -45.0055541992188, 
    -42.591667175293, 
    -48.0444450378418, 
    -35.3583335876465, 
    21.158332824707, 
    23.6499996185303, 
    132.800003051758, 
    381.591674804688, 
    428.433349609375, 
    483.416656494141, 
    624.597229003906, 
    674.116638183594, 
    782.530578613281, 
    969.191650390625, 
    970.875, 
    693.894470214844, 
    739.549987792969, 
    688.191650390625, 
    783.797241210938, 
    193.805160522461, 
    458.25, 
    431.894439697266, 
    131.880508422852, 
    -119.3330078125, 
    -190.661773681641, 
    -250.57926940918, 
    -316.789642333984, 
    -644.506225585938, 
    -1661.10656738281, 
    -2204.29125976562,
  
    -2900.14282226562, 
    -2955.66625976562, 
    -2731.810546875, 
    -2696.458984375, 
    -2671.79541015625, 
    -2652.46704101562, 
    -2723.9130859375, 
    -2616.51049804688, 
    -2537.51318359375, 
    -2550.20336914062, 
    -2511.7705078125, 
    -2509.07153320312, 
    -2327.27563476562, 
    -2052.12719726562, 
    -1816.09741210938, 
    -1964.35913085938, 
    -1923.29748535156, 
    -1721.75341796875, 
    -1802.52954101562, 
    -1980.81091308594, 
    -1658.08190917969, 
    -1603.56591796875, 
    -1533.13903808594, 
    -333.132629394531, 
    -261.118225097656, 
    -253.949493408203, 
    -290.822265625, 
    -382.856201171875, 
    -327.088989257812, 
    -316.625701904297, 
    -297.363128662109, 
    -223.954986572266, 
    -148.364990234375, 
    -35.9087066650391, 
    19.6741714477539, 
    -10.0469236373901, 
    553.422180175781, 
    790.797241210938, 
    696.758361816406, 
    523.744445800781, 
    419.144439697266, 
    363.475006103516, 
    339.072235107422, 
    366.041656494141, 
    339.369445800781, 
    457.29443359375, 
    191.430557250977, 
    63.5888900756836, 
    100.777778625488, 
    207.533340454102, 
    179.894439697266, 
    140.449996948242, 
    79.9250030517578, 
    70.2972259521484, 
    46.6722221374512, 
    -27.6638889312744, 
    20.7250003814697, 
    31.5055561065674, 
    -13.0305557250977, 
    -73.0166702270508, 
    32.1166687011719, 
    37.6444435119629, 
    10.2388887405396, 
    -22.6000003814697, 
    -49.2249984741211, 
    -48.5750007629395, 
    34.0472221374512, 
    131.636108398438, 
    132.127777099609, 
    70.8833312988281, 
    -85.6055526733398, 
    -119.622222900391, 
    -38.9583320617676, 
    33.7333335876465, 
    65.3527755737305, 
    136.522216796875, 
    96.2972259521484, 
    84.6638870239258, 
    172.047225952148, 
    91.8944473266602, 
    9.66388893127441, 
    -37.5444450378418, 
    -124.188888549805, 
    -204.233337402344, 
    -125.349998474121, 
    -99.0888900756836, 
    -65.5527801513672, 
    -78.783332824707, 
    -44.3638877868652, 
    -105.280555725098, 
    -114.75, 
    -92.8305587768555, 
    -70.1555557250977, 
    -60.7555541992188, 
    -59.9111099243164, 
    -78.6500015258789, 
    -69.4388885498047, 
    -15.1333332061768, 
    -36.0472221374512, 
    -103.074996948242, 
    -160.552780151367, 
    -183.125, 
    -145.647216796875, 
    -94.8527755737305, 
    -139.311111450195, 
    -201.875, 
    -120.886108398438, 
    38.9944458007812, 
    -112.758331298828, 
    -8.88055515289307, 
    -29.5861110687256, 
    -84.1416702270508, 
    16.0472221374512, 
    13.5888891220093, 
    24.9333343505859, 
    78.3222198486328, 
    76.9749984741211, 
    71.7972259521484, 
    144.194442749023, 
    255.919448852539, 
    355.825012207031, 
    559.888916015625, 
    658.913879394531, 
    598.188903808594, 
    793.530578613281, 
    854.691650390625, 
    831.04443359375, 
    639.283325195312, 
    321.850006103516, 
    330.285186767578, 
    507.600006103516, 
    901.591674804688, 
    283.183013916016, 
    264.621978759766, 
    2.7743091583252, 
    -132.384368896484, 
    -201.730590820312, 
    -307.598266601562, 
    -761.610473632812, 
    -1766.48449707031, 
    -2140.66748046875,
  
    -2984.39794921875, 
    -2916.5732421875, 
    -2822.13232421875, 
    -2775.04296875, 
    -2750.03100585938, 
    -2756.94604492188, 
    -2818.74780273438, 
    -2729.26489257812, 
    -2658.63232421875, 
    -2665.09130859375, 
    -2590.88427734375, 
    -2475.20361328125, 
    -2358.990234375, 
    -2186.92651367188, 
    -2070.21557617188, 
    -2084.72192382812, 
    -1899.49963378906, 
    -1898.95642089844, 
    -2138.31225585938, 
    -2019.52136230469, 
    -1967.40490722656, 
    -1979.56127929688, 
    -1762.48034667969, 
    -1133.66015625, 
    -223.792953491211, 
    -225.697341918945, 
    -260.6337890625, 
    -325.142578125, 
    -448.6728515625, 
    -570.351440429688, 
    -500.744689941406, 
    -329.130615234375, 
    -258.839691162109, 
    -172.986709594727, 
    -53.5840682983398, 
    8.75394439697266, 
    469.541687011719, 
    1011.67224121094, 
    920.922241210938, 
    721.436096191406, 
    427.819458007812, 
    336.738891601562, 
    427.488891601562, 
    517.6611328125, 
    605.758361816406, 
    380.944458007812, 
    249.405548095703, 
    107.547225952148, 
    120.213890075684, 
    164.616668701172, 
    301.369445800781, 
    353.238891601562, 
    162.777770996094, 
    125.830558776855, 
    107.688888549805, 
    113.041664123535, 
    39.5444450378418, 
    47.0194435119629, 
    113.611106872559, 
    72.0583343505859, 
    38.125, 
    32.8277778625488, 
    14.3222227096558, 
    -19.4861106872559, 
    -31.591667175293, 
    -19.5861110687256, 
    3.0583336353302, 
    105.538887023926, 
    104.85277557373, 
    27.5944442749023, 
    -115.244445800781, 
    -128, 
    -29.6777763366699, 
    90.6444473266602, 
    179.136108398438, 
    213.655548095703, 
    136.024993896484, 
    156.463882446289, 
    174.08610534668, 
    151.727783203125, 
    -26.7250003814697, 
    -92.7111129760742, 
    -111.511108398438, 
    -26.7000007629395, 
    143.588882446289, 
    -19.7749996185303, 
    -98.0083312988281, 
    -60.8833312988281, 
    -40.7361106872559, 
    -8.81388854980469, 
    -113.366668701172, 
    -203.111114501953, 
    -98.1999969482422, 
    -90.3555526733398, 
    -8.53611087799072, 
    1.86944448947906, 
    2.93055558204651, 
    33.658332824707, 
    43.6333351135254, 
    -14.7527780532837, 
    -120.847221374512, 
    -130.908325195312, 
    -121.375, 
    -116.594444274902, 
    -126.25, 
    -80.7277755737305, 
    -49.1500015258789, 
    -38.6749992370605, 
    -115.174995422363, 
    -43.7777786254883, 
    -56.2416648864746, 
    -85.2638854980469, 
    -35.1944427490234, 
    22.5444450378418, 
    44.033332824707, 
    182.58332824707, 
    262.563903808594, 
    205.719451904297, 
    166.572219848633, 
    298.055572509766, 
    509.161102294922, 
    588.927795410156, 
    655.155578613281, 
    728.724975585938, 
    786.849975585938, 
    813.072204589844, 
    739.019470214844, 
    550.399963378906, 
    679.11669921875, 
    951.047241210938, 
    788.691650390625, 
    452.58056640625, 
    346.894439697266, 
    297.223083496094, 
    245.994445800781, 
    -73.4859848022461, 
    -156.841293334961, 
    -253.0263671875, 
    -617.874572753906, 
    -1476.16442871094, 
    -1939.00366210938,
  
    -2937.53198242188, 
    -2916.89135742188, 
    -2947.39916992188, 
    -2883.51049804688, 
    -2846.95239257812, 
    -2866.2841796875, 
    -2863.52685546875, 
    -2815.41772460938, 
    -2786.74926757812, 
    -2723.25390625, 
    -2624.21362304688, 
    -2511.31323242188, 
    -2400.47485351562, 
    -2274.86010742188, 
    -2219.90893554688, 
    -2177.2607421875, 
    -2078.44995117188, 
    -2185.99072265625, 
    -2281.44604492188, 
    -2175.41381835938, 
    -2027.07751464844, 
    -1851.92138671875, 
    -1692.92077636719, 
    -1102.68054199219, 
    -245.987258911133, 
    -228.437927246094, 
    -259.867279052734, 
    -348.7412109375, 
    -478.834991455078, 
    -476.423370361328, 
    -698.468017578125, 
    -651.986511230469, 
    -352.840026855469, 
    -243.89892578125, 
    -141.546005249023, 
    -18.2095050811768, 
    387.508331298828, 
    1069.77221679688, 
    1038.45275878906, 
    974.033325195312, 
    76.4388809204102, 
    488.208343505859, 
    653.7138671875, 
    806.316650390625, 
    882.102783203125, 
    700.397216796875, 
    308.247222900391, 
    71.1222229003906, 
    223.258331298828, 
    459.352783203125, 
    383.950012207031, 
    396.100006103516, 
    186.013885498047, 
    158.969451904297, 
    233.338882446289, 
    222.763885498047, 
    135.438888549805, 
    197.444442749023, 
    175.050003051758, 
    74.8361129760742, 
    23.0499992370605, 
    19.2694454193115, 
    -10.3361110687256, 
    -21.375, 
    -2.65277791023254, 
    10.1138887405396, 
    84.0055541992188, 
    125.427772521973, 
    76.886116027832, 
    -44.8833312988281, 
    -114.155555725098, 
    -50.7305564880371, 
    -71.1083374023438, 
    179.813888549805, 
    227.638885498047, 
    212.272232055664, 
    209.719451904297, 
    122.083335876465, 
    152.930557250977, 
    132.991668701172, 
    31.1777782440186, 
    -48.25, 
    -91.0944442749023, 
    -50.8083343505859, 
    70.4805603027344, 
    26.9444446563721, 
    -64.5611114501953, 
    -49.1638870239258, 
    -133.822219848633, 
    -12.5583333969116, 
    -109.324996948242, 
    -181.505554199219, 
    -32.5166664123535, 
    41.8972244262695, 
    62.8611106872559, 
    77.533332824707, 
    62.6416664123535, 
    98.6972274780273, 
    71.8805541992188, 
    -22.0138893127441, 
    -60.1749992370605, 
    -87.3000030517578, 
    -106.674995422363, 
    -105.988891601562, 
    -68.2388916015625, 
    -15.3249998092651, 
    -23.8861122131348, 
    -54.5250015258789, 
    -55.9722213745117, 
    37.9833335876465, 
    16.6638889312744, 
    1.25833344459534, 
    -14.4805555343628, 
    -1.40277779102325, 
    -6.14166641235352, 
    175.616668701172, 
    284.644439697266, 
    350.497222900391, 
    402.122222900391, 
    261.216674804688, 
    392.897216796875, 
    536.155578613281, 
    744.030578613281, 
    715.433349609375, 
    678.672241210938, 
    720.622192382812, 
    1098.71948242188, 
    649.694458007812, 
    840.20556640625, 
    1214.01391601562, 
    1184.40002441406, 
    966.436096191406, 
    515.25, 
    602.891662597656, 
    552.094421386719, 
    163.052795410156, 
    -108.999374389648, 
    -204.109649658203, 
    -329.999755859375, 
    -973.672607421875, 
    -1745.60400390625,
  
    -2974.9453125, 
    -2964.61547851562, 
    -2958.71313476562, 
    -2956.875, 
    -2942.74731445312, 
    -2929.78100585938, 
    -2902.63916015625, 
    -2875.74926757812, 
    -2822.72583007812, 
    -2744.86450195312, 
    -2674.4033203125, 
    -2584.0625, 
    -2468.27319335938, 
    -2404.43359375, 
    -2388.140625, 
    -2296.6513671875, 
    -2303.29370117188, 
    -2383.921875, 
    -2214.19677734375, 
    -2197.32641601562, 
    -2071.4541015625, 
    -1874.54760742188, 
    -1748.1416015625, 
    -1265.75891113281, 
    -226.397842407227, 
    -220.075546264648, 
    -269.869262695312, 
    -393.521270751953, 
    -696.626831054688, 
    -674.300537109375, 
    -634.192504882812, 
    -560.976196289062, 
    -726.838928222656, 
    -390.127258300781, 
    -232.801727294922, 
    -141.618667602539, 
    271.170867919922, 
    75.4296875, 
    604.6611328125, 
    769.775024414062, 
    360.518463134766, 
    1244.20556640625, 
    1174.73608398438, 
    1106.26110839844, 
    1254.51940917969, 
    1227.2138671875, 
    828.066650390625, 
    577.369445800781, 
    527.222229003906, 
    387.188873291016, 
    391.411102294922, 
    274.508331298828, 
    214.175003051758, 
    308.758331298828, 
    321.41943359375, 
    287.466674804688, 
    250.872222900391, 
    267.563873291016, 
    212.763885498047, 
    86.1777801513672, 
    16.2361106872559, 
    51.4138870239258, 
    43.7666664123535, 
    11.8222217559814, 
    11.6305551528931, 
    97.158332824707, 
    94.2861099243164, 
    118.858329772949, 
    127.125, 
    66.8916625976562, 
    84.3138885498047, 
    57.8277778625488, 
    -9.75, 
    192.29167175293, 
    191.697219848633, 
    222.691665649414, 
    265.394439697266, 
    88.0500030517578, 
    126.466667175293, 
    152.197219848633, 
    37.341667175293, 
    184.891662597656, 
    208.977783203125, 
    69.7083282470703, 
    -90.4583358764648, 
    -51.4583320617676, 
    -57.5833320617676, 
    77.5944442749023, 
    -36.5722236633301, 
    -30.1083335876465, 
    -197.127777099609, 
    -153.727783203125, 
    -53.538890838623, 
    132.558334350586, 
    115.858329772949, 
    104.238891601562, 
    99.1861114501953, 
    149.474990844727, 
    126.833335876465, 
    56.25, 
    24.2555561065674, 
    -35.2027778625488, 
    -95.1222229003906, 
    -118.747222900391, 
    -119.905555725098, 
    -95.4305572509766, 
    -32.6305541992188, 
    -34.3722229003906, 
    -17.2027778625488, 
    45.7249984741211, 
    30.1222229003906, 
    7.87222242355347, 
    -27.3805561065674, 
    -21.5249996185303, 
    57.4916687011719, 
    102.527778625488, 
    149.569442749023, 
    198.855560302734, 
    192.524993896484, 
    119.205558776855, 
    342.430541992188, 
    633.650024414062, 
    544.430541992188, 
    586.805541992188, 
    729.936096191406, 
    1002.12219238281, 
    929.247253417969, 
    559.019470214844, 
    578.327758789062, 
    753.674987792969, 
    670.725036621094, 
    646.005554199219, 
    619.863891601562, 
    412.475006103516, 
    891.116638183594, 
    436.496551513672, 
    -100.980445861816, 
    -152.9970703125, 
    -227.650665283203, 
    -472.357666015625, 
    -940.798400878906,
  
    -3058.96459960938, 
    -3039.125, 
    -3019.17260742188, 
    -2997.96850585938, 
    -2989.3818359375, 
    -2935.91918945312, 
    -2891.92065429688, 
    -2878.67309570312, 
    -2823.5625, 
    -2765.7138671875, 
    -2739.31372070312, 
    -2644.1904296875, 
    -2561.37426757812, 
    -2543.43530273438, 
    -2497.43676757812, 
    -2476.04956054688, 
    -2440.62573242188, 
    -2386.998046875, 
    -2215.73706054688, 
    -2185.66186523438, 
    -2121.3466796875, 
    -1969.40454101562, 
    -1711.20886230469, 
    -1483.47424316406, 
    -235.279373168945, 
    -261.269165039062, 
    -341.097473144531, 
    -400.569061279297, 
    -698.217956542969, 
    -805.379516601562, 
    -448.489166259766, 
    -384.378479003906, 
    -492.631774902344, 
    -335.751403808594, 
    -373.934326171875, 
    -206.460479736328, 
    438.272216796875, 
    270.660705566406, 
    220.206008911133, 
    6.97884559631348, 
    816.586120605469, 
    1412.7666015625, 
    1719.68603515625, 
    1487.43884277344, 
    1670.23327636719, 
    1840.93603515625, 
    1434.45556640625, 
    955.941650390625, 
    401.991668701172, 
    471.952789306641, 
    549.647216796875, 
    495.649993896484, 
    379.916656494141, 
    387.772216796875, 
    361.841674804688, 
    378.372222900391, 
    446.488891601562, 
    399.902770996094, 
    296.377777099609, 
    112.722221374512, 
    -12.9944448471069, 
    138.96110534668, 
    199.891662597656, 
    32.5277786254883, 
    56.9555549621582, 
    74.1388854980469, 
    172.769439697266, 
    144.152786254883, 
    158.722229003906, 
    185.366668701172, 
    8.64166641235352, 
    224.055557250977, 
    188.727783203125, 
    383.011108398438, 
    372.600006103516, 
    310.391662597656, 
    319.397216796875, 
    233.944442749023, 
    152.569442749023, 
    123.963890075684, 
    177.580551147461, 
    216.561111450195, 
    230.655563354492, 
    42.0638885498047, 
    -67.4361114501953, 
    -71.7750015258789, 
    23.6916675567627, 
    -19.8722229003906, 
    -51.086109161377, 
    -107.152778625488, 
    -201.041656494141, 
    -125.313888549805, 
    -70.1666641235352, 
    110.027778625488, 
    97.7666625976562, 
    62.8472213745117, 
    149.113891601562, 
    137.216659545898, 
    140.405548095703, 
    42.6416664123535, 
    70.4416656494141, 
    32.5444450378418, 
    -90.4861068725586, 
    -141.866668701172, 
    -135.280548095703, 
    -85.9972229003906, 
    -168.188888549805, 
    -98.7916641235352, 
    27.8638877868652, 
    47.3611106872559, 
    10.2944440841675, 
    -20.0750007629395, 
    22.4694442749023, 
    37.7972221374512, 
    28.8999996185303, 
    159.96110534668, 
    150.880554199219, 
    91.125, 
    143.050003051758, 
    105.697219848633, 
    243.566665649414, 
    625.061096191406, 
    526.700012207031, 
    815.952758789062, 
    756.069458007812, 
    829.533325195312, 
    652.49169921875, 
    728.488891601562, 
    647.438903808594, 
    913.305541992188, 
    968.75830078125, 
    810.697204589844, 
    398.988891601562, 
    277.105560302734, 
    850.730529785156, 
    682.838928222656, 
    -101.595085144043, 
    -140.106033325195, 
    -194.477645874023, 
    -363.069671630859, 
    -724.30078125,
  
    -3034.47680664062, 
    -3076.55493164062, 
    -3030.90747070312, 
    -3000.37353515625, 
    -2996.66479492188, 
    -2972.33056640625, 
    -2928.78442382812, 
    -2898.06372070312, 
    -2877.61401367188, 
    -2818.037109375, 
    -2774.0146484375, 
    -2724.869140625, 
    -2657.4345703125, 
    -2589.1416015625, 
    -2593.64697265625, 
    -2493.28002929688, 
    -2492.1162109375, 
    -2352.7890625, 
    -2212.3671875, 
    -2083.064453125, 
    -1970.62158203125, 
    -1842.64733886719, 
    -1762.99816894531, 
    -1566.77758789062, 
    -526.893981933594, 
    -278.942474365234, 
    -362.891357421875, 
    -439.319885253906, 
    -570.9775390625, 
    -440.857269287109, 
    -439.687377929688, 
    -351.897674560547, 
    -238.097930908203, 
    -193.239608764648, 
    -211.976577758789, 
    -257.98388671875, 
    26.5848808288574, 
    536.333312988281, 
    902.327758789062, 
    862.680603027344, 
    1045.37219238281, 
    1686.58056640625, 
    1971.28051757812, 
    1607.98059082031, 
    1514.11108398438, 
    1990.80004882812, 
    1734.87780761719, 
    1396.89440917969, 
    1101.26110839844, 
    924.627807617188, 
    786.719421386719, 
    665.650024414062, 
    426.491668701172, 
    357.983337402344, 
    334.344451904297, 
    411.922210693359, 
    528.572204589844, 
    485.644439697266, 
    271.613891601562, 
    164.261108398438, 
    26.5638885498047, 
    160.330551147461, 
    244.733337402344, 
    245.869445800781, 
    145.725006103516, 
    125.969444274902, 
    250.530548095703, 
    265.738891601562, 
    212.96110534668, 
    169.513885498047, 
    89.216667175293, 
    257.311126708984, 
    564.722229003906, 
    582.233337402344, 
    582.461120605469, 
    485.238891601562, 
    384.049987792969, 
    330.555541992188, 
    285.024993896484, 
    346.627777099609, 
    424.394439697266, 
    92.5805587768555, 
    236.113891601562, 
    -39.5222206115723, 
    34.8111114501953, 
    -36.0111122131348, 
    78.4416656494141, 
    -12.4111108779907, 
    -43.4722213745117, 
    63.0055541992188, 
    -61.158332824707, 
    -96.341667175293, 
    -27.1444435119629, 
    126.216667175293, 
    105.847221374512, 
    177.266662597656, 
    248.96110534668, 
    176.630554199219, 
    171.391662597656, 
    155.608337402344, 
    81.5805511474609, 
    138.697219848633, 
    32.211109161377, 
    -166.052780151367, 
    -186.969436645508, 
    -116.27222442627, 
    -69.4388885498047, 
    -7.21388864517212, 
    54.2000007629395, 
    55.2861099243164, 
    30.3500003814697, 
    20.1388893127441, 
    39.5527763366699, 
    52.4527778625488, 
    67.841667175293, 
    167.872222900391, 
    165.688888549805, 
    151.938888549805, 
    183.405548095703, 
    171.322219848633, 
    182.797225952148, 
    372.155548095703, 
    571.3388671875, 
    821.627807617188, 
    575.936096191406, 
    789.236083984375, 
    633.144470214844, 
    367.638885498047, 
    284.380554199219, 
    850.005554199219, 
    815.072204589844, 
    757.541687011719, 
    280.673400878906, 
    442.2861328125, 
    1100.99450683594, 
    786.811096191406, 
    -88.544303894043, 
    -153.051773071289, 
    -242.694427490234, 
    -413.442535400391, 
    -639.620178222656,
  
    -3072.99340820312, 
    -3063.1630859375, 
    -3037.28125, 
    -3025.29321289062, 
    -2996.96948242188, 
    -2978.90087890625, 
    -2934.86474609375, 
    -2904.82153320312, 
    -2888.90551757812, 
    -2867.6669921875, 
    -2808.00610351562, 
    -2750.49340820312, 
    -2721.36303710938, 
    -2635.88549804688, 
    -2611.10424804688, 
    -2525.19604492188, 
    -2501.98876953125, 
    -2371.2841796875, 
    -2215.33837890625, 
    -2153.13134765625, 
    -2102.89331054688, 
    -2024.16650390625, 
    -1963.83386230469, 
    -1873.09655761719, 
    -1654.0732421875, 
    -523.519348144531, 
    -366.487701416016, 
    -413.185882568359, 
    -456.887420654297, 
    -289.603454589844, 
    -470.340484619141, 
    -485.238433837891, 
    -262.054046630859, 
    -198.326232910156, 
    -186.649291992188, 
    -99.601806640625, 
    49.5876350402832, 
    160.100006103516, 
    729.00830078125, 
    1056.59448242188, 
    847.691650390625, 
    1294.61669921875, 
    1696.23889160156, 
    2485.59448242188, 
    2146.76123046875, 
    2171.78051757812, 
    1877.13610839844, 
    1521.34997558594, 
    1408.21118164062, 
    1301.89721679688, 
    990.680541992188, 
    1043.197265625, 
    665.361145019531, 
    235.96110534668, 
    185.552780151367, 
    526.674987792969, 
    746.399963378906, 
    711.5, 
    554.61669921875, 
    341.888885498047, 
    227.705551147461, 
    231.841659545898, 
    249.363891601562, 
    252.980560302734, 
    158.644439697266, 
    165.736114501953, 
    172.936111450195, 
    213.563888549805, 
    299.174987792969, 
    252.436111450195, 
    221.175003051758, 
    476.369445800781, 
    314.222229003906, 
    587.38330078125, 
    749.799987792969, 
    660.072204589844, 
    542.105529785156, 
    528.247253417969, 
    638.427795410156, 
    780.652770996094, 
    566.783325195312, 
    579.063903808594, 
    418.477783203125, 
    391.102783203125, 
    272.713897705078, 
    212.680557250977, 
    262.863891601562, 
    94.3861083984375, 
    195.850006103516, 
    362.672210693359, 
    191.66943359375, 
    107.080558776855, 
    148.408325195312, 
    229.33332824707, 
    180.486114501953, 
    107.025001525879, 
    220.194442749023, 
    223.211120605469, 
    185.108337402344, 
    209.405563354492, 
    174.830551147461, 
    141.261108398438, 
    -46.0249977111816, 
    -156.286117553711, 
    -246.947235107422, 
    -121.819442749023, 
    -47.0055541992188, 
    22.036111831665, 
    60.8666648864746, 
    37.9861106872559, 
    39.1416664123535, 
    61.4861106872559, 
    73.3666687011719, 
    64.4277801513672, 
    109.655555725098, 
    189.716659545898, 
    205.338882446289, 
    258.069458007812, 
    281.433319091797, 
    324.063903808594, 
    373.452789306641, 
    157.058334350586, 
    185.991668701172, 
    214.744445800781, 
    198.630554199219, 
    152.832275390625, 
    468.338623046875, 
    929.305541992188, 
    501.033325195312, 
    769.408325195312, 
    700.4111328125, 
    1105.29443359375, 
    976.966674804688, 
    36.8982887268066, 
    572.066650390625, 
    596.022216796875, 
    -40.3916130065918, 
    -168.384979248047, 
    -277.46923828125, 
    -687.878234863281, 
    -805.0390625,
  
    -3005.82836914062, 
    -2985.27514648438, 
    -2995.13232421875, 
    -2870.69921875, 
    -2899.61279296875, 
    -2969.17041015625, 
    -2939.2216796875, 
    -2900.03271484375, 
    -2879.68530273438, 
    -2835.28247070312, 
    -2820.33618164062, 
    -2758.24975585938, 
    -2721.072265625, 
    -2695.05517578125, 
    -2681.07055664062, 
    -2656.37255859375, 
    -2539.57568359375, 
    -2458.18994140625, 
    -2406.54321289062, 
    -2390.75048828125, 
    -2392.54760742188, 
    -2395.39697265625, 
    -2278.8193359375, 
    -2122.54760742188, 
    -1758.43664550781, 
    -1548.92236328125, 
    -338.316223144531, 
    -385.155944824219, 
    -394.16748046875, 
    -302.926849365234, 
    -462.165130615234, 
    -599.45263671875, 
    -389.096069335938, 
    -245.527954101562, 
    -196.90901184082, 
    -222.82942199707, 
    -108.183792114258, 
    43.9790458679199, 
    184.936111450195, 
    1132.83337402344, 
    1395.19445800781, 
    1139.33605957031, 
    1630.43615722656, 
    2444.52783203125, 
    2392.41674804688, 
    2391.17504882812, 
    1996.4638671875, 
    1479.75830078125, 
    2100.177734375, 
    1794.38610839844, 
    1222.67785644531, 
    1317.47216796875, 
    601.66943359375, 
    225.79167175293, 
    457.769439697266, 
    842.8388671875, 
    1080.31665039062, 
    966.194458007812, 
    860.255554199219, 
    619.805541992188, 
    352.327758789062, 
    324.408325195312, 
    244.844451904297, 
    354.16943359375, 
    228.727783203125, 
    168.352767944336, 
    206.050003051758, 
    288.675018310547, 
    301.54443359375, 
    277.136108398438, 
    146.125, 
    277.977783203125, 
    428.122222900391, 
    468.336120605469, 
    709.086120605469, 
    765.238891601562, 
    855.924987792969, 
    909.108337402344, 
    866.947204589844, 
    665.472229003906, 
    396.20556640625, 
    610.724975585938, 
    793.805541992188, 
    795.375, 
    690.08056640625, 
    258.049987792969, 
    288.833343505859, 
    314.055541992188, 
    485.111114501953, 
    460.072235107422, 
    375.899993896484, 
    206.594451904297, 
    226.980560302734, 
    178.863891601562, 
    89.363883972168, 
    14.9527778625488, 
    67.0222244262695, 
    95.9722213745117, 
    97.1333312988281, 
    190.122222900391, 
    198.686111450195, 
    250.522216796875, 
    127.933326721191, 
    -6.33888912200928, 
    -136.772216796875, 
    -283.219451904297, 
    -112.236114501953, 
    4.71111106872559, 
    18.5722217559814, 
    16.1083335876465, 
    49.6722221374512, 
    87.5055541992188, 
    207.863891601562, 
    155.108337402344, 
    166.027770996094, 
    226.194442749023, 
    292.366668701172, 
    322.047241210938, 
    382.91943359375, 
    486.905548095703, 
    485.91943359375, 
    361.858337402344, 
    75.4694442749023, 
    326.358337402344, 
    678.647216796875, 
    796.424987792969, 
    143.445526123047, 
    388.196594238281, 
    293.891662597656, 
    650.813903808594, 
    761.8388671875, 
    956.494445800781, 
    1068.1611328125, 
    760.891662597656, 
    457.805541992188, 
    568.872253417969, 
    -97.5083694458008, 
    -219.519058227539, 
    -331.242492675781, 
    -820.709350585938, 
    -1104.35705566406,
  
    -2977.11889648438, 
    -2895.24682617188, 
    -3022.66723632812, 
    -2998.99047851562, 
    -2970.91357421875, 
    -2981.6962890625, 
    -2946.22729492188, 
    -2916.76831054688, 
    -2898.8193359375, 
    -2846.87939453125, 
    -2821.57763671875, 
    -2759.61840820312, 
    -2774.12426757812, 
    -2698.28735351562, 
    -2705.33862304688, 
    -2693.61254882812, 
    -2629.072265625, 
    -2613.69091796875, 
    -2558.6923828125, 
    -2552.61669921875, 
    -2585.34228515625, 
    -2490.56591796875, 
    -2333.55615234375, 
    -2116.12182617188, 
    -1826.45166015625, 
    -1812.84362792969, 
    -1356.26733398438, 
    -459.247253417969, 
    -348.69775390625, 
    -309.501190185547, 
    -551.561889648438, 
    -491.290985107422, 
    -190.770843505859, 
    -215.059051513672, 
    -202.216888427734, 
    -278.706024169922, 
    -198.80322265625, 
    -29.7494564056396, 
    457.627655029297, 
    840.244445800781, 
    940.413940429688, 
    1261.06665039062, 
    1840.45275878906, 
    2057.66650390625, 
    2252.26953125, 
    2126.29150390625, 
    1942.4111328125, 
    1731.83056640625, 
    2014.64721679688, 
    2105.86938476562, 
    1603.98889160156, 
    1271.41662597656, 
    1227.67504882812, 
    889.194458007812, 
    1090.13610839844, 
    1163.23889160156, 
    866.702758789062, 
    750.819458007812, 
    968.261108398438, 
    804.066650390625, 
    678.75, 
    432.644439697266, 
    365.075012207031, 
    414.913879394531, 
    337.183319091797, 
    322.808319091797, 
    374.199981689453, 
    357.641662597656, 
    331.563873291016, 
    315.758331298828, 
    264.272216796875, 
    275.447235107422, 
    403.122222900391, 
    559.525024414062, 
    651.730529785156, 
    622.6611328125, 
    865.375, 
    1170.63891601562, 
    986.905578613281, 
    790.086120605469, 
    752.9638671875, 
    716.030578613281, 
    606.858337402344, 
    425.16943359375, 
    67.9472198486328, 
    116.675003051758, 
    133.530548095703, 
    378.75, 
    462.258331298828, 
    528.652770996094, 
    474.252777099609, 
    433.325012207031, 
    409.027770996094, 
    359.699981689453, 
    110.541664123535, 
    2.64166641235352, 
    89.4749984741211, 
    -8.19444465637207, 
    161.300003051758, 
    151.772216796875, 
    207.725006103516, 
    349.030548095703, 
    272.375, 
    181.138885498047, 
    -4.38611030578613, 
    -166.502777099609, 
    -73.1444473266602, 
    -27.2972221374512, 
    -37.9638900756836, 
    -17.1333332061768, 
    122.997222900391, 
    178.16667175293, 
    240.766662597656, 
    226.147216796875, 
    240.797225952148, 
    293.438873291016, 
    331.375, 
    383.555541992188, 
    441.244445800781, 
    560.194458007812, 
    652.54443359375, 
    589.166625976562, 
    261.519439697266, 
    711.119445800781, 
    906.827819824219, 
    689.197204589844, 
    485.933319091797, 
    -48.4356498718262, 
    192.179122924805, 
    693, 
    748.033325195312, 
    940.174987792969, 
    1156.54443359375, 
    320.438873291016, 
    419.522216796875, 
    696.355529785156, 
    -101.638000488281, 
    -242.654067993164, 
    -327.650054931641, 
    -660.636840820312, 
    -981.414733886719,
  
    -2922.23095703125, 
    -2837.67724609375, 
    -2872.42309570312, 
    -2972.83935546875, 
    -2988.61767578125, 
    -2980.21044921875, 
    -2933.32543945312, 
    -2916.32958984375, 
    -2904.02490234375, 
    -2854.04125976562, 
    -2835.87084960938, 
    -2794.82739257812, 
    -2774.1787109375, 
    -2776.05639648438, 
    -2751.04296875, 
    -2740.75366210938, 
    -2743.09106445312, 
    -2678.88500976562, 
    -2620.3505859375, 
    -2613.6318359375, 
    -2632.09399414062, 
    -2512.1220703125, 
    -2388.3916015625, 
    -2231.10107421875, 
    -2120.4560546875, 
    -2038.69445800781, 
    -1836.2939453125, 
    -1531.02429199219, 
    -513.418212890625, 
    -354.295501708984, 
    -557.361389160156, 
    -383.754302978516, 
    -224.115005493164, 
    -217.917770385742, 
    -272.819946289062, 
    -277.693298339844, 
    -251.464721679688, 
    -204.300750732422, 
    -113.177680969238, 
    156.569961547852, 
    456.219451904297, 
    1413.87219238281, 
    1539.43334960938, 
    1610.26391601562, 
    2530.03881835938, 
    2292.33325195312, 
    2132.14428710938, 
    1474.09716796875, 
    1498.34448242188, 
    2035.28051757812, 
    1802.68884277344, 
    1662.16943359375, 
    1265.42224121094, 
    873.602783203125, 
    1394.34448242188, 
    1503.84448242188, 
    765.780517578125, 
    868.502746582031, 
    1310.7861328125, 
    1444.96105957031, 
    1007.44720458984, 
    629.816650390625, 
    503.438873291016, 
    479.638885498047, 
    360.824981689453, 
    396.933319091797, 
    382.761108398438, 
    251.438888549805, 
    432.255554199219, 
    448.477783203125, 
    309.149993896484, 
    228.669448852539, 
    311.552795410156, 
    449.899993896484, 
    536.302795410156, 
    499.116668701172, 
    546.011108398438, 
    1052.322265625, 
    784.422241210938, 
    678.486083984375, 
    929.880554199219, 
    842.119445800781, 
    535.238891601562, 
    326.744445800781, 
    657.269470214844, 
    586.238891601562, 
    558.722229003906, 
    515.069458007812, 
    404.611114501953, 
    452.780548095703, 
    553.663879394531, 
    649.188903808594, 
    547.308349609375, 
    360.061126708984, 
    143.988891601562, 
    117.966667175293, 
    352.413879394531, 
    148.680557250977, 
    -53.7111129760742, 
    78.7083358764648, 
    4.67777681350708, 
    236.619445800781, 
    315.019439697266, 
    266.566650390625, 
    263.325012207031, 
    191.655548095703, 
    116.85277557373, 
    21.8333339691162, 
    66.6194458007812, 
    104.805557250977, 
    224.927780151367, 
    215.858337402344, 
    229.716659545898, 
    213.097213745117, 
    231.03889465332, 
    327.461120605469, 
    370.905548095703, 
    420.386108398438, 
    457.844451904297, 
    559.4638671875, 
    762.536071777344, 
    603.25830078125, 
    724.7861328125, 
    76.2611083984375, 
    624.436096191406, 
    843.269409179688, 
    881.291687011719, 
    744.473083496094, 
    -9.40828514099121, 
    673.724975585938, 
    649.174987792969, 
    689.130554199219, 
    778.258361816406, 
    772.269409179688, 
    -72.0247116088867, 
    132.005752563477, 
    -194.473129272461, 
    -534.597045898438, 
    -953.666442871094, 
    -767.976806640625, 
    -907.292785644531,
  
    -2981.2841796875, 
    -2876.11791992188, 
    -2914.13427734375, 
    -2920.39575195312, 
    -2990.43237304688, 
    -2980.7373046875, 
    -2973.93994140625, 
    -2931.951171875, 
    -2916.21948242188, 
    -2881.03637695312, 
    -2883.36181640625, 
    -2853.58813476562, 
    -2814.57177734375, 
    -2809.14404296875, 
    -2805.72583007812, 
    -2829.28686523438, 
    -2768.13671875, 
    -2752.96533203125, 
    -2708.76928710938, 
    -2692.12646484375, 
    -2611.94067382812, 
    -2576.96411132812, 
    -2488.07250976562, 
    -2431.64892578125, 
    -2329.49340820312, 
    -2178.99877929688, 
    -1988.60607910156, 
    -1749.84985351562, 
    -1415.64233398438, 
    -403.387329101562, 
    -385.949523925781, 
    -366.952239990234, 
    -369.523590087891, 
    -258.370849609375, 
    -254.422836303711, 
    -296.878204345703, 
    -298.638671875, 
    -278.466522216797, 
    -313.265258789062, 
    -288.150848388672, 
    395.620086669922, 
    911.4111328125, 
    1262.58605957031, 
    1658.4638671875, 
    2081.57495117188, 
    2252.58056640625, 
    2094.25830078125, 
    1693.74719238281, 
    1345.27783203125, 
    2025.52502441406, 
    2052.9638671875, 
    1951.26391601562, 
    1558.55554199219, 
    1535.65002441406, 
    1298.09729003906, 
    1227.30004882812, 
    706.158325195312, 
    1234.91662597656, 
    1287.22497558594, 
    1165.24169921875, 
    945.172241210938, 
    677.63330078125, 
    604.311157226562, 
    548.974975585938, 
    489.913879394531, 
    391.108337402344, 
    424.369445800781, 
    409.447204589844, 
    427.716674804688, 
    549.041687011719, 
    425.608337402344, 
    337.072204589844, 
    282.558349609375, 
    399.605560302734, 
    734.977783203125, 
    542.627807617188, 
    621.763854980469, 
    818.79443359375, 
    853.002807617188, 
    1058.55004882812, 
    1216.61669921875, 
    1208.14453125, 
    813.327758789062, 
    615.41943359375, 
    1115.16662597656, 
    1008.75830078125, 
    835.255554199219, 
    761.150024414062, 
    382.269439697266, 
    376.961120605469, 
    595.238891601562, 
    573.299987792969, 
    409.941680908203, 
    279.969451904297, 
    166.194442749023, 
    208.547225952148, 
    237.425003051758, 
    219.644439697266, 
    73.1194458007812, 
    -16.4499988555908, 
    268.538879394531, 
    19.125, 
    290.066650390625, 
    333.569458007812, 
    304.508331298828, 
    261.113891601562, 
    243.20832824707, 
    88.8916702270508, 
    -94.6222229003906, 
    116.29167175293, 
    112.261108398438, 
    145.736114501953, 
    138.588882446289, 
    145.497222900391, 
    202.269439697266, 
    339.297210693359, 
    416.336120605469, 
    469.902770996094, 
    664.716674804688, 
    621.591674804688, 
    826.875, 
    704.416625976562, 
    810.333374023438, 
    726.308349609375, 
    -76.2111206054688, 
    506.752777099609, 
    721.288879394531, 
    789.116638183594, 
    -48.2354774475098, 
    550, 
    547.297241210938, 
    477.944427490234, 
    300.263885498047, 
    650.969482421875, 
    190.726119995117, 
    -176.617767333984, 
    -365.656524658203, 
    -1062.78173828125, 
    -2495.49829101562, 
    -2889.181640625, 
    -2235.7939453125,
  
    -3067.703125, 
    -2798.3984375, 
    -2765.4091796875, 
    -2965.6474609375, 
    -2985.68041992188, 
    -2755.03759765625, 
    -2955.50366210938, 
    -2917.37060546875, 
    -2936.82666015625, 
    -2901.7119140625, 
    -2891.43530273438, 
    -2876.265625, 
    -2879.86669921875, 
    -2920.27734375, 
    -2836.79248046875, 
    -2837.81982421875, 
    -2786.62963867188, 
    -2777.34497070312, 
    -2782.35400390625, 
    -2689.0908203125, 
    -2685.65405273438, 
    -2603.61254882812, 
    -2596.32250976562, 
    -2499.28881835938, 
    -2393.1923828125, 
    -2280.24658203125, 
    -2077.92553710938, 
    -1826.09631347656, 
    -1702.09509277344, 
    -1389.86279296875, 
    -1013.76159667969, 
    -1064.17272949219, 
    -693.096313476562, 
    -309.613037109375, 
    -267.871215820312, 
    -321.421783447266, 
    -272.485626220703, 
    -283.623413085938, 
    -258.550811767578, 
    -194.926727294922, 
    -88.3203277587891, 
    195.591674804688, 
    823.858337402344, 
    1212.47497558594, 
    1595.26940917969, 
    1666.61669921875, 
    1659.99169921875, 
    1546.32775878906, 
    1727.55834960938, 
    1746.75561523438, 
    1825.9638671875, 
    1814.86389160156, 
    1776.36108398438, 
    1685.86389160156, 
    942.597229003906, 
    969.658325195312, 
    1060.26940917969, 
    1379.96948242188, 
    1222.63061523438, 
    1092.69165039062, 
    799.552795410156, 
    647.377746582031, 
    658.5361328125, 
    638.95556640625, 
    616.813903808594, 
    568.091674804688, 
    522.049987792969, 
    606.716674804688, 
    592.933349609375, 
    520.172241210938, 
    458.030548095703, 
    375.416656494141, 
    318.813903808594, 
    319.191680908203, 
    470.794464111328, 
    507.072235107422, 
    727.569458007812, 
    946.902770996094, 
    1113.33325195312, 
    1248.64440917969, 
    1313.86389160156, 
    1170.7861328125, 
    1173.19165039062, 
    992.277770996094, 
    1174.84167480469, 
    1008.38610839844, 
    743.952758789062, 
    475.111114501953, 
    392.436096191406, 
    413.269439697266, 
    602.022216796875, 
    526.108337402344, 
    491.936126708984, 
    401.022216796875, 
    333.5, 
    405.355560302734, 
    245.366668701172, 
    276.488891601562, 
    77.7138900756836, 
    -166.752777099609, 
    -116.602783203125, 
    174.227783203125, 
    264.311126708984, 
    241.04167175293, 
    259.197235107422, 
    324.005554199219, 
    302.350006103516, 
    258.138885498047, 
    257.452758789062, 
    71.9305572509766, 
    106.683334350586, 
    83.1611099243164, 
    111.616668701172, 
    165.477783203125, 
    140.280548095703, 
    344.613891601562, 
    446.788909912109, 
    499.024993896484, 
    585.380554199219, 
    706.252746582031, 
    696.813903808594, 
    920.563903808594, 
    566.7138671875, 
    641.722229003906, 
    415.188873291016, 
    72.7436981201172, 
    418.808349609375, 
    481.811126708984, 
    -40.5645408630371, 
    443.394439697266, 
    428.663879394531, 
    391.605560302734, 
    489.050018310547, 
    19.5130424499512, 
    -142.921188354492, 
    -322.499877929688, 
    -847.838012695312, 
    -1309.9794921875, 
    -2142.01953125, 
    -2168.31640625, 
    -1615.49560546875,
  
    -3108.58178710938, 
    -2879.13647460938, 
    -2830.4384765625, 
    -3004.71362304688, 
    -3006.64306640625, 
    -2969.19311523438, 
    -2965.56811523438, 
    -2876.97216796875, 
    -2951.3017578125, 
    -2923.64624023438, 
    -2910.66577148438, 
    -2884.2109375, 
    -2872.1611328125, 
    -2895.07348632812, 
    -2889.1650390625, 
    -2806.46875, 
    -2797.3798828125, 
    -2780.64331054688, 
    -2774.28051757812, 
    -2717.97802734375, 
    -2677.46630859375, 
    -2648.99072265625, 
    -2614.11010742188, 
    -2565.5361328125, 
    -2445.74731445312, 
    -2319.20654296875, 
    -2150.64233398438, 
    -1941.43994140625, 
    -1868.55712890625, 
    -1670.28576660156, 
    -1410.1328125, 
    -1139.28295898438, 
    -831.148132324219, 
    -316.854736328125, 
    -249.530883789062, 
    -267.026245117188, 
    -338.444854736328, 
    -245.715194702148, 
    -289.304107666016, 
    -276.027374267578, 
    -284.941589355469, 
    -164.528350830078, 
    -10.04660987854, 
    386.673309326172, 
    702.469421386719, 
    836.549987792969, 
    1034.95275878906, 
    1083.20837402344, 
    1269.55834960938, 
    1650.75280761719, 
    1853.95556640625, 
    1308.822265625, 
    1464.69995117188, 
    1182.26953125, 
    646.772216796875, 
    904.663879394531, 
    847.755554199219, 
    1034.03332519531, 
    1079.322265625, 
    1043.65551757812, 
    813.825012207031, 
    763.0361328125, 
    749.08056640625, 
    708.88330078125, 
    778.791687011719, 
    787.058349609375, 
    524.79443359375, 
    563.372253417969, 
    619.741638183594, 
    579.147216796875, 
    538.136108398438, 
    548.105529785156, 
    421.622222900391, 
    335.772216796875, 
    403.174987792969, 
    492.647216796875, 
    690.561096191406, 
    877.983337402344, 
    1022.74444580078, 
    1103.00561523438, 
    1268.94165039062, 
    1396.10278320312, 
    1104.677734375, 
    790.847229003906, 
    760.863891601562, 
    594.9638671875, 
    763.519409179688, 
    689.061096191406, 
    546.219421386719, 
    442.480560302734, 
    501.600006103516, 
    470.200012207031, 
    365.052764892578, 
    422.924987792969, 
    434.811126708984, 
    299.450012207031, 
    444.591674804688, 
    451.391662597656, 
    237.83610534668, 
    214.399993896484, 
    10.2972230911255, 
    -159.366668701172, 
    212.66667175293, 
    30.1749992370605, 
    184.369445800781, 
    172.102783203125, 
    255.675003051758, 
    193.21110534668, 
    283.738891601562, 
    122.436111450195, 
    206, 
    156.933334350586, 
    42.25, 
    96.7972183227539, 
    34.3916664123535, 
    212.322219848633, 
    354.116668701172, 
    489.405548095703, 
    438.322204589844, 
    250.433334350586, 
    472.827789306641, 
    547.849975585938, 
    455.022216796875, 
    734.930541992188, 
    672.766662597656, 
    387.219451904297, 
    -11.233775138855, 
    139.370559692383, 
    -46.4845733642578, 
    106.554000854492, 
    283.061126708984, 
    215.711120605469, 
    325.413879394531, 
    56.413028717041, 
    -292.807891845703, 
    -1288.27819824219, 
    -1941.02185058594, 
    -2051.65966796875, 
    -2197.111328125, 
    -2279.51147460938, 
    -3280.19360351562,
  
    -2954.32934570312, 
    -2858.318359375, 
    -3090.6728515625, 
    -3098.74780273438, 
    -2928.07690429688, 
    -2965.310546875, 
    -2899.19018554688, 
    -2911.42846679688, 
    -2940.34814453125, 
    -2880.94091796875, 
    -2912.45751953125, 
    -2892.97387695312, 
    -2879.93603515625, 
    -2875.13647460938, 
    -2848.6123046875, 
    -2877.60107421875, 
    -2815.03466796875, 
    -2789.5126953125, 
    -2775.69921875, 
    -2766.82153320312, 
    -2725.29931640625, 
    -2693.19702148438, 
    -2693.5400390625, 
    -2610.6396484375, 
    -2517.4091796875, 
    -2407.27563476562, 
    -2340.72216796875, 
    -2147.09497070312, 
    -2009.95300292969, 
    -1754.28845214844, 
    -1483.82250976562, 
    -1163.650390625, 
    -945.311645507812, 
    -640.09375, 
    -252.400405883789, 
    -213.950576782227, 
    -267.773376464844, 
    -302.81396484375, 
    -301.786346435547, 
    -306.315460205078, 
    -339.894317626953, 
    -241.818603515625, 
    -190.392776489258, 
    -148.942657470703, 
    -60.3312873840332, 
    241.704025268555, 
    95.6472244262695, 
    410.372222900391, 
    780.288879394531, 
    1365.01391601562, 
    1679.53332519531, 
    1645.27221679688, 
    1588.302734375, 
    1058.69165039062, 
    413.575012207031, 
    713.041625976562, 
    1520.72497558594, 
    1463.18054199219, 
    1210.65270996094, 
    999.677795410156, 
    953.819458007812, 
    911.736145019531, 
    952.572204589844, 
    868.130554199219, 
    935.594421386719, 
    893.75, 
    689.913879394531, 
    642.052795410156, 
    646.600036621094, 
    650.405517578125, 
    523.833312988281, 
    711.086120605469, 
    817.563903808594, 
    940.683349609375, 
    524.136108398438, 
    480.583343505859, 
    947.549987792969, 
    913.280517578125, 
    999.447204589844, 
    944.511108398438, 
    1412.7138671875, 
    1395.13330078125, 
    1350.23327636719, 
    1120.20275878906, 
    907.844421386719, 
    1015.46667480469, 
    1202.75830078125, 
    966.524963378906, 
    840.7138671875, 
    561.666687011719, 
    512.163879394531, 
    712.79443359375, 
    632.147216796875, 
    661.488891601562, 
    613.333312988281, 
    418.583343505859, 
    452.680541992188, 
    445.822204589844, 
    460.352783203125, 
    215.805557250977, 
    321.66943359375, 
    94.1888885498047, 
    150.636108398438, 
    294.816680908203, 
    372.138885498047, 
    293.788879394531, 
    342.58056640625, 
    146.347229003906, 
    208.966659545898, 
    114.222221374512, 
    63.783332824707, 
    11.4388885498047, 
    8.34166622161865, 
    -50.9972229003906, 
    -62.6833305358887, 
    116.108329772949, 
    308.702789306641, 
    338.030548095703, 
    256.758331298828, 
    325.522216796875, 
    327.975006103516, 
    316.538879394531, 
    703.552734375, 
    848.052795410156, 
    340.666656494141, 
    660.066650390625, 
    402.352783203125, 
    19.5635833740234, 
    68.2053527832031, 
    -79.3710479736328, 
    88.6920928955078, 
    171.319442749023, 
    284.530548095703, 
    -58.468334197998, 
    -185.878616333008, 
    -1550.14050292969, 
    -3049.95556640625, 
    -3162.14575195312, 
    -3054.70239257812, 
    -3468.04907226562, 
    -3603.73779296875,
  
    -2851.56201171875, 
    -2551.37280273438, 
    -2766.728515625, 
    -2986.64013671875, 
    -2806.19409179688, 
    -2989.52270507812, 
    -2725.82885742188, 
    -2915.79052734375, 
    -2915.857421875, 
    -2714.31298828125, 
    -2899.17333984375, 
    -2893.8037109375, 
    -2902.36083984375, 
    -2893.72875976562, 
    -2891.6552734375, 
    -2867.63745117188, 
    -2863.244140625, 
    -2827.2265625, 
    -2803.70336914062, 
    -2786.95947265625, 
    -2775.24169921875, 
    -2742.77587890625, 
    -2726.37768554688, 
    -2706.96264648438, 
    -2648.58862304688, 
    -2550.64575195312, 
    -2454.01513671875, 
    -2304.2255859375, 
    -2104.84814453125, 
    -1883.78698730469, 
    -1608.67578125, 
    -1375.80993652344, 
    -1302.54565429688, 
    -1023.28466796875, 
    -553.270385742188, 
    -290.219635009766, 
    -275.157684326172, 
    -298.975067138672, 
    -299.472259521484, 
    -303.552337646484, 
    -308.770660400391, 
    -294.063079833984, 
    -284.527313232422, 
    -283.717407226562, 
    -254.508255004883, 
    -198.748291015625, 
    -142.647857666016, 
    -70.2449951171875, 
    280.859741210938, 
    811.555541992188, 
    1040.47216796875, 
    1021.31109619141, 
    1245.38610839844, 
    273.374206542969, 
    1370.72216796875, 
    2105.26928710938, 
    2226.74731445312, 
    1903.21948242188, 
    1549.49169921875, 
    1363.23327636719, 
    1278.48889160156, 
    1280.33056640625, 
    1140.32495117188, 
    1143.48059082031, 
    1075.36108398438, 
    969.019470214844, 
    840.494445800781, 
    755.672241210938, 
    698.650024414062, 
    665.38330078125, 
    642.033325195312, 
    564.805541992188, 
    1051.83325195312, 
    1196.77770996094, 
    1099.41943359375, 
    620.702758789062, 
    987.569458007812, 
    1170.59448242188, 
    1496.05834960938, 
    1552.66943359375, 
    1642.13610839844, 
    1829.78063964844, 
    1731.95275878906, 
    1532.93896484375, 
    1526.32495117188, 
    1488.98059082031, 
    1223.27502441406, 
    1281.32495117188, 
    1044.08605957031, 
    622.36669921875, 
    405.875, 
    684.638916015625, 
    803.877807617188, 
    856.4111328125, 
    715.255554199219, 
    648.566650390625, 
    519.900024414062, 
    621.577758789062, 
    626.49169921875, 
    342.047210693359, 
    415.352752685547, 
    464.758331298828, 
    130.202774047852, 
    311.513885498047, 
    177.652770996094, 
    221.205551147461, 
    6.9611120223999, 
    -91.4833374023438, 
    84.6611099243164, 
    -28.7194442749023, 
    278.613891601562, 
    -115.511116027832, 
    -181.133331298828, 
    -220.297225952148, 
    -107.697219848633, 
    -16.1833324432373, 
    62.0388870239258, 
    -12.2138891220093, 
    337.197235107422, 
    182.761108398438, 
    71.783332824707, 
    353.575012207031, 
    718.299987792969, 
    281.5, 
    232.436111450195, 
    564.894470214844, 
    624.166687011719, 
    193.608337402344, 
    237.786117553711, 
    -70.33203125, 
    -96.206901550293, 
    -27.2295837402344, 
    32.0001068115234, 
    -101.972579956055, 
    -127.035980224609, 
    -507.338256835938, 
    -3022.87255859375, 
    -3260.611328125, 
    -3335.02221679688, 
    -3535.26416015625, 
    -3613.6953125,
  
    -2899.98559570312, 
    -2451.96362304688, 
    -2661.33251953125, 
    -2492.5693359375, 
    -2690.75927734375, 
    -2870.80810546875, 
    -2935.2138671875, 
    -2625.08325195312, 
    -2986.32080078125, 
    -2909.65795898438, 
    -2942.95678710938, 
    -2876.5615234375, 
    -2837.1025390625, 
    -2898.9794921875, 
    -2889.98266601562, 
    -2889.21533203125, 
    -2866.53442382812, 
    -2847.23876953125, 
    -2863.86010742188, 
    -2899.55541992188, 
    -2811.55517578125, 
    -2782.34204101562, 
    -2787.37182617188, 
    -2736.60034179688, 
    -2705.7861328125, 
    -2645.45239257812, 
    -2542.11743164062, 
    -2385.34594726562, 
    -2218.9794921875, 
    -2065.2392578125, 
    -1807.65283203125, 
    -1639.2880859375, 
    -1604.84509277344, 
    -1441.79650878906, 
    -1111.18176269531, 
    -458.014404296875, 
    -259.865936279297, 
    -282.868499755859, 
    -292.935485839844, 
    -298.108581542969, 
    -298.825714111328, 
    -342.083404541016, 
    -316.86572265625, 
    -353.320770263672, 
    -390.160583496094, 
    -298.587829589844, 
    -184.607070922852, 
    -150.468521118164, 
    -93.1434173583984, 
    4.07357788085938, 
    655.650024414062, 
    172.808334350586, 
    162.637084960938, 
    1077.93884277344, 
    1944.40551757812, 
    2123.86108398438, 
    2365.16943359375, 
    2346.51391601562, 
    1974.56945800781, 
    1333.66394042969, 
    1457.12780761719, 
    1422.427734375, 
    1486.39721679688, 
    1431.68615722656, 
    1265.33618164062, 
    1085.47229003906, 
    1004.18609619141, 
    1093.77502441406, 
    1032.96118164062, 
    816.594482421875, 
    953.997253417969, 
    1088.14440917969, 
    1201.2861328125, 
    1180.22497558594, 
    1297.78332519531, 
    1191.93054199219, 
    1276.06945800781, 
    1216.15283203125, 
    1462.46105957031, 
    1375.04162597656, 
    1791.61950683594, 
    2041.59448242188, 
    1874.34997558594, 
    1523.76672363281, 
    1855.05554199219, 
    1633.17224121094, 
    1470.52770996094, 
    1415.22778320312, 
    1042.85278320312, 
    941.266662597656, 
    726.7861328125, 
    790.966674804688, 
    797.941650390625, 
    1071.95556640625, 
    761.869445800781, 
    758.772216796875, 
    683.799987792969, 
    884.125, 
    970.288879394531, 
    244.047225952148, 
    618.572204589844, 
    546.441650390625, 
    286.877777099609, 
    102.29167175293, 
    220.486114501953, 
    155.183334350586, 
    307.102783203125, 
    -127.549995422363, 
    -162.816665649414, 
    -284.941650390625, 
    -249.33332824707, 
    -288.924987792969, 
    -203.572219848633, 
    -151.919448852539, 
    -30.3166656494141, 
    103.130554199219, 
    126.586112976074, 
    275.011108398438, 
    462.408325195312, 
    464.725006103516, 
    517.9111328125, 
    372.241668701172, 
    259.490264892578, 
    9.27665233612061, 
    12.4472055435181, 
    192.734115600586, 
    303.666717529297, 
    17.2383117675781, 
    -89.5387573242188, 
    -126.92008972168, 
    -124.836334228516, 
    -108.115211486816, 
    -103.248497009277, 
    -90.7778701782227, 
    -111.843284606934, 
    -385.016326904297, 
    -2093.70385742188, 
    -2562.11865234375, 
    -3303.08081054688, 
    -3591.1611328125, 
    -3698.55517578125,
  
    -2828.48876953125, 
    -2652.58056640625, 
    -2677.6640625, 
    -2563.32397460938, 
    -2648.53442382812, 
    -2839.544921875, 
    -2870.67553710938, 
    -2847.99853515625, 
    -2981.25, 
    -2834.62817382812, 
    -2902.4755859375, 
    -2872.544921875, 
    -2805.771484375, 
    -2874.95556640625, 
    -2891.68920898438, 
    -2798.61401367188, 
    -2872.81274414062, 
    -2854.11669921875, 
    -2833.51708984375, 
    -2863.0810546875, 
    -2867.61767578125, 
    -2780.92724609375, 
    -2806.68969726562, 
    -2770.2138671875, 
    -2747.62231445312, 
    -2710.36669921875, 
    -2645.61352539062, 
    -2460.06225585938, 
    -2350.40991210938, 
    -2161.93969726562, 
    -2001.73474121094, 
    -1923.69946289062, 
    -1785.77014160156, 
    -1683.11340332031, 
    -1463.04541015625, 
    -890.018432617188, 
    -299.082794189453, 
    -324.717895507812, 
    -279.011779785156, 
    -285.752746582031, 
    -297.589447021484, 
    -305.391448974609, 
    -324.177764892578, 
    -393.535461425781, 
    -358.356079101562, 
    -208.292221069336, 
    -201.260299682617, 
    -196.198822021484, 
    -235.699188232422, 
    -251.928359985352, 
    -425.462921142578, 
    537.566345214844, 
    1213.48608398438, 
    1384.12219238281, 
    1852.25830078125, 
    2129.29443359375, 
    2297.43603515625, 
    2474.80541992188, 
    2158.79711914062, 
    1911.21667480469, 
    1783.40002441406, 
    1142.31945800781, 
    1609.052734375, 
    1579.69995117188, 
    1468.26940917969, 
    1323.61938476562, 
    1138.67224121094, 
    1404.5361328125, 
    1493.2666015625, 
    1211.53051757812, 
    1037.35827636719, 
    1314.77502441406, 
    1799.16662597656, 
    1480.40270996094, 
    1566.01672363281, 
    1432.99450683594, 
    1434.25830078125, 
    1339.55004882812, 
    1125.66943359375, 
    1830.70275878906, 
    2074.78881835938, 
    1924.75561523438, 
    1960.63891601562, 
    2128.0166015625, 
    1977.70556640625, 
    1610.11669921875, 
    1527.29174804688, 
    1569.77221679688, 
    1487.09716796875, 
    1320.85559082031, 
    984.844421386719, 
    835.927795410156, 
    943.04443359375, 
    1137.01672363281, 
    936.66943359375, 
    764.980529785156, 
    745.388854980469, 
    1121.13330078125, 
    1064.17492675781, 
    786.530517578125, 
    1064.23327636719, 
    985.030578613281, 
    463.744445800781, 
    249.502777099609, 
    426.261108398438, 
    532.527770996094, 
    276.186096191406, 
    72.5527801513672, 
    -180.655563354492, 
    -275.222229003906, 
    -305.338897705078, 
    -374.436126708984, 
    -325.16943359375, 
    -234.377777099609, 
    -51.7999992370605, 
    110.902778625488, 
    300.491668701172, 
    523.191650390625, 
    259.647216796875, 
    623.958312988281, 
    681.522216796875, 
    904.58056640625, 
    891.563903808594, 
    675.255554199219, 
    578.238891601562, 
    198.463470458984, 
    84.6900177001953, 
    16.5818309783936, 
    -78.9966049194336, 
    27.5252590179443, 
    -105.035308837891, 
    -107.410697937012, 
    -101.457252502441, 
    -101.267372131348, 
    -125.948394775391, 
    -848.986083984375, 
    -2277.76904296875, 
    -2592.3876953125, 
    -3599.19677734375, 
    -2481.01196289062, 
    -3389.49072265625,
  
    -2481.46948242188, 
    -2428.31372070312, 
    -2701.5810546875, 
    -2822.21118164062, 
    -2531.59814453125, 
    -2740.20092773438, 
    -2661.94897460938, 
    -2708.22387695312, 
    -2856.1875, 
    -2700.90991210938, 
    -2736.9892578125, 
    -2613.98999023438, 
    -2738.025390625, 
    -2702.97241210938, 
    -2894.15161132812, 
    -2872.71850585938, 
    -2896.3623046875, 
    -2887.119140625, 
    -2890.13745117188, 
    -2830.78125, 
    -2852.3193359375, 
    -2795.78735351562, 
    -2814.00048828125, 
    -2807.53247070312, 
    -2805.16381835938, 
    -2741.50317382812, 
    -2693.1875, 
    -2594.90698242188, 
    -2515.82104492188, 
    -2360.60595703125, 
    -2223.98217773438, 
    -2156.720703125, 
    -2033.99633789062, 
    -1890.39611816406, 
    -1608.59350585938, 
    -1190.41540527344, 
    -596.234619140625, 
    -272.995941162109, 
    -279.1142578125, 
    -279.683929443359, 
    -291.807830810547, 
    -300.406311035156, 
    -300.709045410156, 
    -329.0615234375, 
    -278.148071289062, 
    -256.200439453125, 
    -314.754547119141, 
    -394.9482421875, 
    -440.67626953125, 
    -460.330688476562, 
    -229.447219848633, 
    299.561096191406, 
    915.147216796875, 
    1392.2333984375, 
    1750.75280761719, 
    2033.15002441406, 
    2401.62768554688, 
    2352.13623046875, 
    2260.7138671875, 
    2355.06103515625, 
    2085.31665039062, 
    1576.81665039062, 
    1392.05554199219, 
    1305.5888671875, 
    1588.97497558594, 
    1473.25549316406, 
    915.819458007812, 
    1299.802734375, 
    1750.15551757812, 
    1773.77502441406, 
    922.313903808594, 
    1301.96667480469, 
    1411.2861328125, 
    1316.69165039062, 
    1503.52502441406, 
    1110.06945800781, 
    1648.3583984375, 
    1632.32495117188, 
    1767.48608398438, 
    1878.84448242188, 
    1746.85559082031, 
    1503.86389160156, 
    1677.12219238281, 
    1741.20007324219, 
    1809.63049316406, 
    1791.99719238281, 
    1258.81115722656, 
    1468.20556640625, 
    1360.87219238281, 
    1071.1416015625, 
    888.741638183594, 
    919.002746582031, 
    957.525024414062, 
    785.133361816406, 
    878.358337402344, 
    850.9638671875, 
    1506.62219238281, 
    1805.93054199219, 
    1525.36389160156, 
    875.113891601562, 
    1213.61938476562, 
    1273.86389160156, 
    646.58056640625, 
    252.808334350586, 
    75.6555557250977, 
    163.449996948242, 
    278.144439697266, 
    480.980560302734, 
    327.222229003906, 
    74.0861129760742, 
    68.1638870239258, 
    -76.6194381713867, 
    -255.752777099609, 
    -224.972213745117, 
    -228.96110534668, 
    -29.3638896942139, 
    224.572219848633, 
    488.233337402344, 
    800.458312988281, 
    147.055557250977, 
    405.733337402344, 
    209.925003051758, 
    411.438873291016, 
    609.527770996094, 
    480.377777099609, 
    408.786102294922, 
    110.81364440918, 
    0.737175166606903, 
    -1.24231207370758, 
    -5.60969877243042, 
    -142.157028198242, 
    -125.415687561035, 
    -146.350952148438, 
    -256.174011230469, 
    -825.412170410156, 
    -2673.0703125, 
    -2834.77807617188, 
    -3382.65502929688, 
    -3535.54956054688, 
    -3617.64965820312, 
    -4006.548828125,
  
    -2476.47241210938, 
    -2352.85620117188, 
    -2368.90063476562, 
    -2417.92651367188, 
    -2386.42358398438, 
    -2436.80346679688, 
    -2433.81103515625, 
    -2473.56567382812, 
    -2592.56103515625, 
    -2649.77661132812, 
    -2558.97485351562, 
    -2659.03466796875, 
    -2548.37622070312, 
    -2702.70288085938, 
    -2804.0517578125, 
    -2650.962890625, 
    -2671.82958984375, 
    -2652.20043945312, 
    -2891.54638671875, 
    -2885.21459960938, 
    -2604.00903320312, 
    -2811.2998046875, 
    -2813.27978515625, 
    -2815.62451171875, 
    -2812.45434570312, 
    -2763.39038085938, 
    -2712.40307617188, 
    -2668.02880859375, 
    -2611.619140625, 
    -2478.34838867188, 
    -2394.05322265625, 
    -2304.29565429688, 
    -2188.96142578125, 
    -1995.87280273438, 
    -1608.71081542969, 
    -1190.51159667969, 
    -630.708190917969, 
    -298.054901123047, 
    -320.115936279297, 
    -328.259124755859, 
    -321.517272949219, 
    -311.263671875, 
    -374.098510742188, 
    -389.723846435547, 
    -324.357147216797, 
    -391.722595214844, 
    -561.1630859375, 
    -515.254516601562, 
    -491.321868896484, 
    -389.934020996094, 
    -175.450225830078, 
    536.611083984375, 
    355.513885498047, 
    1153.46667480469, 
    314.644439697266, 
    590.836120605469, 
    1416.09448242188, 
    1863.47778320312, 
    1842.01940917969, 
    2319.34155273438, 
    2363.322265625, 
    1947.09448242188, 
    1755.51391601562, 
    1393.99719238281, 
    1176.15551757812, 
    1649.61389160156, 
    1771.61389160156, 
    1232.43884277344, 
    1735.09716796875, 
    1611.66943359375, 
    1456.63610839844, 
    1244.17785644531, 
    1400.95007324219, 
    1396.88049316406, 
    1570.98889160156, 
    1546.93054199219, 
    1496.40832519531, 
    1488.65002441406, 
    2216.40551757812, 
    1846.20556640625, 
    1712.35278320312, 
    1742.2861328125, 
    2003.88049316406, 
    1477.13891601562, 
    1524.50280761719, 
    1707.27783203125, 
    1645.05554199219, 
    1500.13061523438, 
    677.799987792969, 
    1304.04443359375, 
    764.813903808594, 
    670.866638183594, 
    855.972229003906, 
    1216.75280761719, 
    1350.66394042969, 
    1619.98608398438, 
    1603.93615722656, 
    1659.0888671875, 
    1830.625, 
    1718.947265625, 
    1213.85827636719, 
    1409.99169921875, 
    1201.64721679688, 
    859.944458007812, 
    434.494445800781, 
    394.644439697266, 
    810.969421386719, 
    675.75, 
    775.716674804688, 
    688.688903808594, 
    835.802795410156, 
    361.763885498047, 
    -75.5611114501953, 
    -315.205535888672, 
    -124.66389465332, 
    -304.447235107422, 
    46.1527786254883, 
    667.150024414062, 
    561.461120605469, 
    390.327789306641, 
    897.611083984375, 
    879.341674804688, 
    318.980560302734, 
    920.155578613281, 
    456.602783203125, 
    394.333312988281, 
    175.563888549805, 
    -1.58709251880646, 
    -43.2000885009766, 
    -104.091171264648, 
    -117.84252166748, 
    -131.293228149414, 
    -205.592910766602, 
    -1332.44982910156, 
    -2506.34936523438, 
    -2945.00341796875, 
    -3281.53735351562, 
    -3342.8203125, 
    -3482.54370117188, 
    -3905.62841796875, 
    -3859.29931640625,
  
    -2329.44311523438, 
    -2250.97778320312, 
    -2336.64526367188, 
    -2407.8515625, 
    -2391.29028320312, 
    -2389.28588867188, 
    -2436.55297851562, 
    -2387.95703125, 
    -2556.75512695312, 
    -2567.39013671875, 
    -2366.11767578125, 
    -2508.56127929688, 
    -2545.30224609375, 
    -2695.57641601562, 
    -2633.45263671875, 
    -2538.14184570312, 
    -2508.12744140625, 
    -2620.017578125, 
    -2712.13500976562, 
    -2793.91162109375, 
    -2803.7470703125, 
    -2633.4775390625, 
    -2779.46166992188, 
    -2811.05883789062, 
    -2795.0419921875, 
    -2747.22802734375, 
    -2709.85034179688, 
    -2709.50024414062, 
    -2650.62255859375, 
    -2572.25903320312, 
    -2498.021484375, 
    -2410.00659179688, 
    -2293.4326171875, 
    -2085.7509765625, 
    -1580.44140625, 
    -1148.21923828125, 
    -486.322845458984, 
    -345.794372558594, 
    -400.819488525391, 
    -425.743499755859, 
    -474.123382568359, 
    -467.645416259766, 
    -483.827819824219, 
    -500.704223632812, 
    -508.365844726562, 
    -622.991149902344, 
    -597.519836425781, 
    -431.872497558594, 
    -376.923217773438, 
    -306.706848144531, 
    -198.39501953125, 
    60.2056465148926, 
    236.136108398438, 
    -118.716667175293, 
    974, 
    1601.42504882812, 
    1828.375, 
    1671.15283203125, 
    2030.11669921875, 
    2303.55541992188, 
    2381.15283203125, 
    2313.24169921875, 
    1769.02221679688, 
    1053.98608398438, 
    1327.89440917969, 
    1325.1611328125, 
    1149.09997558594, 
    554.363891601562, 
    1450.81115722656, 
    1270.75561523438, 
    1203.34729003906, 
    1610, 
    1217.7333984375, 
    505.106048583984, 
    1681.65551757812, 
    1749.35278320312, 
    1357.17504882812, 
    1141.23059082031, 
    1704.38342285156, 
    1796.24719238281, 
    1415.78894042969, 
    1415.34448242188, 
    1514.0166015625, 
    1073.95275878906, 
    1691.71667480469, 
    1509.75, 
    1473.76672363281, 
    1506.447265625, 
    1373.00549316406, 
    1072.8583984375, 
    897.311096191406, 
    1143.67785644531, 
    995.344421386719, 
    579.094421386719, 
    1343.96948242188, 
    1851.06384277344, 
    1543.18334960938, 
    1368.0361328125, 
    1073.29724121094, 
    1407.70556640625, 
    1053.96105957031, 
    878.2861328125, 
    671.111083984375, 
    621.29443359375, 
    73.3472213745117, 
    362.736114501953, 
    729.766662597656, 
    629.349975585938, 
    265.950012207031, 
    162.241668701172, 
    526.005554199219, 
    453.255554199219, 
    -286.733337402344, 
    -238.111114501953, 
    441.786102294922, 
    677.358337402344, 
    -158.350006103516, 
    -19.7930297851562, 
    107.340812683105, 
    168.166427612305, 
    260.702789306641, 
    867.430541992188, 
    301.933837890625, 
    880.233337402344, 
    776.655578613281, 
    784.122192382812, 
    454.699981689453, 
    349.891662597656, 
    32.62353515625, 
    -54.258975982666, 
    -101.447364807129, 
    -113.175033569336, 
    -203.583587646484, 
    -1057.68395996094, 
    -2647.49853515625, 
    -2736.32373046875, 
    -3220.06298828125, 
    -3241.37280273438, 
    -3596.71801757812, 
    -3720.96240234375, 
    -3199.1337890625,
  
    -2300, 
    -2297.22021484375, 
    -2181.25122070312, 
    -2270.66552734375, 
    -2220.49389648438, 
    -2269.8701171875, 
    -2388.3447265625, 
    -2407.31591796875, 
    -2381.99145507812, 
    -2373.95971679688, 
    -2327.62036132812, 
    -2447.28002929688, 
    -2554.97509765625, 
    -2351.41650390625, 
    -2439.49609375, 
    -2565.990234375, 
    -2463.49853515625, 
    -2509.59057617188, 
    -2593.92041015625, 
    -2643.42138671875, 
    -2759.20556640625, 
    -2533.04541015625, 
    -2676.40502929688, 
    -2709.8994140625, 
    -2747.7392578125, 
    -2787.66772460938, 
    -2733.69116210938, 
    -2679.13452148438, 
    -2713.4521484375, 
    -2615.06518554688, 
    -2533.810546875, 
    -2460.04541015625, 
    -2301.1572265625, 
    -2068.80981445312, 
    -1567.86779785156, 
    -1101.33068847656, 
    -498.89599609375, 
    -397.627075195312, 
    -423.793884277344, 
    -458.706085205078, 
    -492.733215332031, 
    -444.692169189453, 
    -439.055755615234, 
    -433.47314453125, 
    -425.226165771484, 
    -387.0830078125, 
    -241.098648071289, 
    -163.094024658203, 
    -241.545303344727, 
    -295.507507324219, 
    -258.686950683594, 
    -165.729904174805, 
    89.8868103027344, 
    405.599975585938, 
    1348.88891601562, 
    1789.375, 
    2219.61401367188, 
    2079.03881835938, 
    2048.74169921875, 
    2477.84448242188, 
    2424.20556640625, 
    1978.16394042969, 
    1370.61389160156, 
    1202.64721679688, 
    901.62841796875, 
    796.552062988281, 
    1544.99719238281, 
    1174.13891601562, 
    1148.34997558594, 
    1360.50280761719, 
    1523.60278320312, 
    931.513916015625, 
    1270.5546875, 
    499.402160644531, 
    1827.96118164062, 
    1623.322265625, 
    1131.45837402344, 
    1373.29162597656, 
    574.900024414062, 
    1509.17736816406, 
    621.540344238281, 
    583.523559570312, 
    1428.93884277344, 
    1793.4111328125, 
    1646.98327636719, 
    1199.70837402344, 
    1444.427734375, 
    1522.88891601562, 
    1730.12219238281, 
    1369.60559082031, 
    1090.38610839844, 
    1338.17492675781, 
    756.08056640625, 
    852.655578613281, 
    1257.90002441406, 
    1248.40832519531, 
    1111.15283203125, 
    1110.89453125, 
    904.736083984375, 
    925.5888671875, 
    676.208312988281, 
    799.349975585938, 
    429.263885498047, 
    19.4055557250977, 
    -236.180557250977, 
    423.100006103516, 
    526.216674804688, 
    408.524993896484, 
    308.355560302734, 
    184.927780151367, 
    30.9333343505859, 
    182.184326171875, 
    -41.3698692321777, 
    -259.347229003906, 
    589.619445800781, 
    461.302795410156, 
    -21.9329509735107, 
    0.783912777900696, 
    529.700012207031, 
    226.492477416992, 
    126.359764099121, 
    346.236114501953, 
    -37.1607551574707, 
    109.794799804688, 
    535.752807617188, 
    670.244445800781, 
    385.744445800781, 
    537.841674804688, 
    284.477783203125, 
    248.485397338867, 
    -174.455352783203, 
    -105.212829589844, 
    -212.967071533203, 
    -1610.19616699219, 
    -2928.82934570312, 
    -3082.32006835938, 
    -3146.96630859375, 
    -3299.03076171875, 
    -3652.37524414062, 
    -2841.94750976562, 
    -2569.88452148438,
  
    -2300, 
    -2292.49780273438, 
    -1982.38244628906, 
    -2096.50170898438, 
    -2217.38037109375, 
    -2242.95361328125, 
    -2325.64794921875, 
    -2174.99389648438, 
    -2231.3505859375, 
    -2358.23046875, 
    -2372.6904296875, 
    -2363.28198242188, 
    -2361.02001953125, 
    -2419.568359375, 
    -2504.34790039062, 
    -2400.45727539062, 
    -2274.43505859375, 
    -2497.50732421875, 
    -2461.75219726562, 
    -2524.46435546875, 
    -2371.32153320312, 
    -2631.69384765625, 
    -2510.64331054688, 
    -2493.33569335938, 
    -2510.4599609375, 
    -2523.26123046875, 
    -2619.91772460938, 
    -2667.11303710938, 
    -2675.2041015625, 
    -2609.90087890625, 
    -2538.60009765625, 
    -2438.14697265625, 
    -2302.37475585938, 
    -2157.86303710938, 
    -1707.94311523438, 
    -1229.03735351562, 
    -554.143127441406, 
    -410.123809814453, 
    -410.791839599609, 
    -418.482421875, 
    -411.80419921875, 
    -398.318695068359, 
    -348.446868896484, 
    -323.901916503906, 
    -305.556182861328, 
    -247.754776000977, 
    -214.449279785156, 
    -181.373443603516, 
    -202.925201416016, 
    -257.218048095703, 
    -303.148162841797, 
    -359.873352050781, 
    29.9130573272705, 
    551.516662597656, 
    954.638854980469, 
    1843.875, 
    1723.46667480469, 
    1994.74169921875, 
    2170.67504882812, 
    2429, 
    2358.533203125, 
    2232.822265625, 
    1353.45556640625, 
    1330.19165039062, 
    1083.92224121094, 
    -234.763427734375, 
    774.287841796875, 
    414.948791503906, 
    583.342956542969, 
    634.808349609375, 
    1048.822265625, 
    845.093627929688, 
    -476.9501953125, 
    2032.28881835938, 
    1553.79162597656, 
    1875.95275878906, 
    1517.80554199219, 
    1707.63891601562, 
    1168.09448242188, 
    1418.28332519531, 
    692.146423339844, 
    754.516357421875, 
    1855.87219238281, 
    1799.9638671875, 
    1275.19995117188, 
    946.502807617188, 
    992.147216796875, 
    1409.99719238281, 
    1622.73608398438, 
    1253.90832519531, 
    1254.95275878906, 
    1223.89172363281, 
    1041.58056640625, 
    1059.49719238281, 
    810.752746582031, 
    595.363891601562, 
    120.405555725098, 
    258.288879394531, 
    75.3249969482422, 
    94.6500015258789, 
    227.483337402344, 
    -241.263885498047, 
    -303.227783203125, 
    -305.455535888672, 
    -77.2555541992188, 
    27.0027770996094, 
    27.3552703857422, 
    11.7891235351562, 
    7.64732122421265, 
    -18.6361198425293, 
    -21.6966934204102, 
    -29.2650356292725, 
    7.99591493606567, 
    -111.100006103516, 
    59.4415588378906, 
    -16.7220096588135, 
    -84.7085571289062, 
    -112.462287902832, 
    403.291625976562, 
    219.002258300781, 
    -127.861938476562, 
    431.258331298828, 
    206.566757202148, 
    202.22721862793, 
    260.766662597656, 
    300.16943359375, 
    310.191650390625, 
    273.336120605469, 
    333.100006103516, 
    181.167098999023, 
    -184.681381225586, 
    -98.4742736816406, 
    -516.123901367188, 
    -2582.40307617188, 
    -2964.0498046875, 
    -3065.41625976562, 
    -3173.04931640625, 
    -3044.10668945312, 
    -3149.85913085938, 
    -3477.54467773438, 
    -3284.34619140625,
  
    -2300, 
    -2300, 
    -2193.22607421875, 
    -1839.00549316406, 
    -1890.23229980469, 
    -2039.59484863281, 
    -2195.51831054688, 
    -2239.1064453125, 
    -2264.44580078125, 
    -2162.94799804688, 
    -2263.80590820312, 
    -2288.09252929688, 
    -2187.94653320312, 
    -2215.92211914062, 
    -2366.908203125, 
    -2404.72314453125, 
    -2360.64379882812, 
    -2228.35034179688, 
    -2329.17749023438, 
    -2319.00048828125, 
    -2307.36059570312, 
    -2523.99340820312, 
    -2366.93579101562, 
    -2392.2509765625, 
    -2399.31298828125, 
    -2403.70581054688, 
    -2418.8955078125, 
    -2410.74951171875, 
    -2499.4580078125, 
    -2492.67895507812, 
    -2438.95825195312, 
    -2389.01049804688, 
    -2319.4560546875, 
    -2224.11206054688, 
    -1860.1640625, 
    -1367.9052734375, 
    -775.429870605469, 
    -366.008544921875, 
    -361.346160888672, 
    -309.984252929688, 
    -292.585296630859, 
    -313.051696777344, 
    -312.367645263672, 
    -305.531890869141, 
    -310.226501464844, 
    -283.521179199219, 
    -263.549713134766, 
    -222.591079711914, 
    -207.976470947266, 
    -245.858779907227, 
    -281.950103759766, 
    -285.986267089844, 
    -203.850555419922, 
    73.7556533813477, 
    1307.69995117188, 
    1131.8388671875, 
    1829.0361328125, 
    1839.18884277344, 
    2306.91381835938, 
    2431.36108398438, 
    2190.36108398438, 
    1891.45837402344, 
    679.408325195312, 
    449.587005615234, 
    1523.57507324219, 
    712.952270507812, 
    780.949401855469, 
    1113.8896484375, 
    1199.61938476562, 
    1677.58056640625, 
    1632.11938476562, 
    -309.950958251953, 
    1043.37219238281, 
    1742.72497558594, 
    1552.01672363281, 
    1915.75, 
    1034.90270996094, 
    1402.38891601562, 
    -235.112777709961, 
    1184.00280761719, 
    924.107116699219, 
    445.402526855469, 
    1394.80554199219, 
    1372.56945800781, 
    644.900024414062, 
    1245.36950683594, 
    280.055541992188, 
    1079.72497558594, 
    1491.49169921875, 
    884.727783203125, 
    802.450012207031, 
    1179.80554199219, 
    1212.78051757812, 
    1299.08337402344, 
    1309.79724121094, 
    585.319458007812, 
    499.630554199219, 
    560.027770996094, 
    342.038909912109, 
    190.630554199219, 
    20.9500980377197, 
    32.0717124938965, 
    248.105560302734, 
    421.186126708984, 
    378.244445800781, 
    401.308319091797, 
    333.761108398438, 
    392.726348876953, 
    -4.16288614273071, 
    -21.8262748718262, 
    -4.98491287231445, 
    -29.5834293365479, 
    0.871506929397583, 
    -29.9629650115967, 
    -78.4756317138672, 
    -93.9791946411133, 
    -177.26188659668, 
    -196.102905273438, 
    -198.824325561523, 
    -182.733779907227, 
    -290.769348144531, 
    -194.440795898438, 
    -109.166435241699, 
    -115.071800231934, 
    -22.5695915222168, 
    -53.5741729736328, 
    146.96110534668, 
    111.438888549805, 
    344.994445800781, 
    -1.30565714836121, 
    -109.526916503906, 
    -435.500915527344, 
    -2270.56298828125, 
    -2807.73193359375, 
    -3019.34057617188, 
    -3217.244140625, 
    -3692.99975585938, 
    -4574.02734375, 
    -3466.35107421875, 
    -3231.38500976562, 
    -2933.55810546875,
  
    -2300, 
    -2300, 
    -2300, 
    -1865.90466308594, 
    -1822.71838378906, 
    -1864.26745605469, 
    -1885.09753417969, 
    -1987.04968261719, 
    -2121.20166015625, 
    -2183.2353515625, 
    -2268.71362304688, 
    -2166.53881835938, 
    -2207.0517578125, 
    -2209.98608398438, 
    -2154.8701171875, 
    -2167.07958984375, 
    -2154.6669921875, 
    -2238.591796875, 
    -2337.63354492188, 
    -2288.23168945312, 
    -2246.88500976562, 
    -2341.17211914062, 
    -2343.77172851562, 
    -2288.69677734375, 
    -2302.7861328125, 
    -2197.15087890625, 
    -2199.3740234375, 
    -2243.40844726562, 
    -2312.01171875, 
    -2288.1796875, 
    -2262.95458984375, 
    -2249.18359375, 
    -2189.76538085938, 
    -2093.48217773438, 
    -1922.47436523438, 
    -1557.5712890625, 
    -1211.82861328125, 
    -573.013366699219, 
    -340.610870361328, 
    -306.498046875, 
    -295.154663085938, 
    -297.977020263672, 
    -310.635375976562, 
    -315.033233642578, 
    -308.155181884766, 
    -296.002471923828, 
    -301.858795166016, 
    -264.453460693359, 
    -263.332397460938, 
    -296.523101806641, 
    -264.170654296875, 
    -281.851623535156, 
    -273.211273193359, 
    -192.591583251953, 
    296.672210693359, 
    808.947204589844, 
    1530.13330078125, 
    1576.9638671875, 
    2568.96655273438, 
    2351.94165039062, 
    2078.81103515625, 
    1919.81396484375, 
    729.091674804688, 
    -636.986450195312, 
    756.361572265625, 
    335.826568603516, 
    1384.2666015625, 
    1333.59167480469, 
    993.900756835938, 
    1640.71105957031, 
    2052.02783203125, 
    29.4036502838135, 
    1518.62219238281, 
    2330.2861328125, 
    666.761108398438, 
    1744.39172363281, 
    1349.30554199219, 
    1233.13330078125, 
    1261.20275878906, 
    119.592979431152, 
    588.961120605469, 
    1300.84997558594, 
    540.837707519531, 
    403.715423583984, 
    738.424987792969, 
    411.138885498047, 
    376.430541992188, 
    716.400024414062, 
    980.752807617188, 
    801.038879394531, 
    1218.65270996094, 
    1469.58056640625, 
    1161.072265625, 
    1599.2666015625, 
    1430.60278320312, 
    847.061096191406, 
    699.119445800781, 
    749.075012207031, 
    534.586120605469, 
    563.630554199219, 
    10.9703969955444, 
    81.6227340698242, 
    460.188903808594, 
    209.486099243164, 
    811.636108398438, 
    188.292633056641, 
    27.8870582580566, 
    167.944442749023, 
    7.30294942855835, 
    25.0968647003174, 
    18.9765930175781, 
    -34.9095306396484, 
    -30.9417667388916, 
    -62.3214416503906, 
    -92.6266784667969, 
    -139.738494873047, 
    -205.231658935547, 
    -200.825271606445, 
    -203.073806762695, 
    -193.941024780273, 
    -174.847839355469, 
    -172.789138793945, 
    -267.635864257812, 
    -260.913269042969, 
    -164.435852050781, 
    -84.7320251464844, 
    -81.8106307983398, 
    -35.1345176696777, 
    -55.3474044799805, 
    -118.504592895508, 
    -159.433944702148, 
    -1242.3271484375, 
    -2908.9384765625, 
    -2914.67553710938, 
    -3174.64672851562, 
    -3347.74780273438, 
    -4386.81689453125, 
    -3274.65356445312, 
    -2731.97729492188, 
    -3624.43603515625, 
    -4296.65283203125,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1712.93957519531, 
    -1710.56555175781, 
    -1747.06970214844, 
    -1817.79833984375, 
    -1801.99328613281, 
    -1856.03295898438, 
    -2024.3740234375, 
    -2242.43188476562, 
    -2244.70239257812, 
    -2141.20581054688, 
    -2122.17431640625, 
    -2088.0380859375, 
    -2112.16186523438, 
    -2067.11010742188, 
    -2111.75024414062, 
    -2198.90014648438, 
    -2296.49145507812, 
    -2169.34619140625, 
    -2078.28125, 
    -2165.37670898438, 
    -2286.7939453125, 
    -2107.93310546875, 
    -2107.6806640625, 
    -2145.18237304688, 
    -2096.1123046875, 
    -1967.34631347656, 
    -1969.92541503906, 
    -1907.43518066406, 
    -1779.54846191406, 
    -1761.16162109375, 
    -1798.54357910156, 
    -1584.82470703125, 
    -1376.24206542969, 
    -1110.70422363281, 
    -848.210754394531, 
    -408.879150390625, 
    -322.989318847656, 
    -294.609313964844, 
    -303.366058349609, 
    -320.294708251953, 
    -310.702087402344, 
    -325.820434570312, 
    -315.205627441406, 
    -288.154876708984, 
    -292.412658691406, 
    -263.161651611328, 
    -268.420684814453, 
    -312.5380859375, 
    -544.922180175781, 
    -264.184936523438, 
    103.276519775391, 
    772.397216796875, 
    1359.55834960938, 
    1621.72216796875, 
    2523.18603515625, 
    2390.591796875, 
    1957.31945800781, 
    1584.11389160156, 
    1004.9638671875, 
    1774.10559082031, 
    528.286865234375, 
    1276.18884277344, 
    1073.25646972656, 
    1890.37219238281, 
    691.834594726562, 
    1297.38720703125, 
    1245.51953125, 
    711.859558105469, 
    1185.9111328125, 
    1997.29443359375, 
    1102.05004882812, 
    659.616638183594, 
    267.216583251953, 
    1155.88330078125, 
    960.850402832031, 
    -92.79541015625, 
    -105.228591918945, 
    777.7861328125, 
    566.350891113281, 
    -128.97119140625, 
    42.2875480651855, 
    632.652770996094, 
    363.272216796875, 
    948.727783203125, 
    439.830535888672, 
    1389.02502441406, 
    1560.56665039062, 
    1334.49438476562, 
    1148.77502441406, 
    1193.46667480469, 
    987.291687011719, 
    445.411346435547, 
    1032.2861328125, 
    335.841674804688, 
    673.002807617188, 
    61.6408920288086, 
    28.8414344787598, 
    -50.5800895690918, 
    6.84631586074829, 
    144.516662597656, 
    263.236114501953, 
    -77.0827789306641, 
    206.476501464844, 
    -19.6784725189209, 
    -68.6207656860352, 
    -111.135932922363, 
    -161.542144775391, 
    -171.575698852539, 
    -216.726379394531, 
    -302.891235351562, 
    -292.288360595703, 
    -156.385665893555, 
    -80.295295715332, 
    -96.5050582885742, 
    -93.0644836425781, 
    -82.7820587158203, 
    -46.7531929016113, 
    -135.240463256836, 
    -181.618255615234, 
    -271.306976318359, 
    -178.826263427734, 
    -119.863784790039, 
    -87.5197067260742, 
    -60.4147148132324, 
    -48.8173332214355, 
    -116.89070892334, 
    -596.368103027344, 
    -2479.69140625, 
    -2860.51147460938, 
    -3150.92553710938, 
    -3386.20922851562, 
    -3996.21850585938, 
    -4312.99951171875, 
    -3074.46264648438, 
    -3200.09252929688, 
    -4147.9951171875, 
    -4383.3935546875,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1654.267578125, 
    -1646.2841796875, 
    -1651.29040527344, 
    -1706.11462402344, 
    -1672.283203125, 
    -1749.54968261719, 
    -1837.08459472656, 
    -1921.22094726562, 
    -2091.68212890625, 
    -2170.43896484375, 
    -2106.76977539062, 
    -2088.09204101562, 
    -2084.35864257812, 
    -1988.73034667969, 
    -1965.86901855469, 
    -2013.119140625, 
    -2009.685546875, 
    -2035.0205078125, 
    -2147.1220703125, 
    -2110.87646484375, 
    -1929.63269042969, 
    -2035.19958496094, 
    -1900.07458496094, 
    -1835.20629882812, 
    -1801.11560058594, 
    -1651.55554199219, 
    -1575.19604492188, 
    -1279.48937988281, 
    -1332.61975097656, 
    -1457.85180664062, 
    -1402.14428710938, 
    -1380.98034667969, 
    -1192.62048339844, 
    -991.917114257812, 
    -593.665283203125, 
    -430.042907714844, 
    -342.639434814453, 
    -331.212554931641, 
    -332.478424072266, 
    -313.280181884766, 
    -339.720001220703, 
    -328.260223388672, 
    -309.753692626953, 
    -301.759643554688, 
    -283.542144775391, 
    -237.62028503418, 
    -342.437133789062, 
    -411.304473876953, 
    -201.239990234375, 
    -173.998718261719, 
    173.595489501953, 
    627.797241210938, 
    1056.65002441406, 
    1600.9111328125, 
    1934.19445800781, 
    1874.84716796875, 
    1575.3388671875, 
    1523.51110839844, 
    1424.64172363281, 
    358.398071289062, 
    -480.882446289062, 
    87.536979675293, 
    893.605529785156, 
    1036.97216796875, 
    28.0311470031738, 
    82.2202072143555, 
    -128.151947021484, 
    1811.85278320312, 
    1607.53051757812, 
    1848.052734375, 
    1618.38330078125, 
    1206.73889160156, 
    -309.128814697266, 
    452.924530029297, 
    1159.13891601562, 
    537.107055664062, 
    722.611083984375, 
    664.906982421875, 
    390.154632568359, 
    317, 
    826.827758789062, 
    679.022216796875, 
    426.002777099609, 
    914.227783203125, 
    1542.18054199219, 
    849.599975585938, 
    1293.24450683594, 
    472.936096191406, 
    995.077819824219, 
    661.842590332031, 
    1070.16943359375, 
    889.049987792969, 
    667.307495117188, 
    708.847229003906, 
    19.9515991210938, 
    -65.8765869140625, 
    -154.419876098633, 
    -13.9557218551636, 
    239.580551147461, 
    350.608337402344, 
    32.5069847106934, 
    -114.051620483398, 
    18.2925910949707, 
    27.2653503417969, 
    -189.429290771484, 
    -301.316741943359, 
    -304.986572265625, 
    -310.066711425781, 
    -258.360046386719, 
    -160.612335205078, 
    -55.5358657836914, 
    -46.51953125, 
    -30.0032501220703, 
    -63.942211151123, 
    -120.341148376465, 
    -178.077255249023, 
    -108.907302856445, 
    -171.762588500977, 
    -158.106552124023, 
    -170.585968017578, 
    -183.539672851562, 
    -161.660827636719, 
    -71.5111083984375, 
    -66.1542663574219, 
    -281.589691162109, 
    -1120.59594726562, 
    -2783.63452148438, 
    -3148.8671875, 
    -3153.63720703125, 
    -3512.96826171875, 
    -4146.1357421875, 
    -3391.62377929688, 
    -2223.818359375, 
    -3364.90112304688, 
    -4007.12133789062, 
    -3707.31298828125,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2280.3095703125, 
    -1523.36157226562, 
    -1544.51538085938, 
    -1684.75671386719, 
    -1663.80187988281, 
    -1693.6025390625, 
    -1736.46704101562, 
    -1682.67565917969, 
    -1768.09265136719, 
    -1886.05847167969, 
    -2042.92565917969, 
    -2076.34033203125, 
    -2002.9921875, 
    -1986.95837402344, 
    -1972.23828125, 
    -1895.03552246094, 
    -1903.654296875, 
    -1889.26354980469, 
    -1999.337890625, 
    -2041.97583007812, 
    -1925.203125, 
    -1835.04382324219, 
    -1824.09912109375, 
    -1683.65502929688, 
    -1601.32666015625, 
    -1526.53601074219, 
    -1378.71789550781, 
    -1295.56396484375, 
    -1255.71594238281, 
    -1219.56066894531, 
    -1179.03112792969, 
    -1178.88830566406, 
    -1034.80480957031, 
    -953.387756347656, 
    -705.70068359375, 
    -497.492095947266, 
    -466.571899414062, 
    -355.765350341797, 
    -367.989196777344, 
    -348.996978759766, 
    -365.246551513672, 
    -349.958679199219, 
    -330.919097900391, 
    -318.300018310547, 
    -270.079162597656, 
    -298.480438232422, 
    -391.005340576172, 
    -254.23649597168, 
    -204.862976074219, 
    -290.495269775391, 
    -170.92204284668, 
    544, 
    1099.21105957031, 
    1561.85278320312, 
    1693.86669921875, 
    1589.18054199219, 
    1470.78332519531, 
    1459.0888671875, 
    1739.21948242188, 
    1493.22497558594, 
    777.544189453125, 
    -598.824523925781, 
    93.3644104003906, 
    -451.717376708984, 
    -409.842498779297, 
    -441.640502929688, 
    222.628890991211, 
    823.091674804688, 
    702.638916015625, 
    1003.78332519531, 
    1044.18884277344, 
    314.653564453125, 
    -296.599060058594, 
    351.958343505859, 
    499.344451904297, 
    759.319458007812, 
    413.010284423828, 
    -261.722991943359, 
    1044.21118164062, 
    814.569396972656, 
    710.525024414062, 
    1195.23059082031, 
    153.314682006836, 
    151.313888549805, 
    516.224975585938, 
    1326.38049316406, 
    900.691650390625, 
    728.014831542969, 
    839.476318359375, 
    862.146545410156, 
    882.147216796875, 
    685.952758789062, 
    707.780517578125, 
    44.7807960510254, 
    -181.492156982422, 
    -182.224685668945, 
    257.919738769531, 
    15.7344102859497, 
    195.688888549805, 
    88.7732467651367, 
    -84.2141647338867, 
    -170.635223388672, 
    -142.769653320312, 
    -132.592010498047, 
    -347.650848388672, 
    -480.272888183594, 
    -375.138824462891, 
    -166.407623291016, 
    -59.4749946594238, 
    -59.9434471130371, 
    -58.7569885253906, 
    -52.9888076782227, 
    -106.175216674805, 
    -151.294097900391, 
    -196.387878417969, 
    -186.33723449707, 
    -138.835647583008, 
    -110.289756774902, 
    -148.712539672852, 
    -168.353485107422, 
    -195.779891967773, 
    -120.839393615723, 
    -62.7992706298828, 
    -231.162887573242, 
    -1529.20007324219, 
    -2534.96240234375, 
    -3060.22875976562, 
    -3221.98608398438, 
    -3747.36474609375, 
    -4018.23315429688, 
    -3700.603515625, 
    -2548.94604492188, 
    -2723.95239257812, 
    -3458.173828125, 
    -2645.44384765625, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2110.1337890625, 
    -1485.87158203125, 
    -1534.44030761719, 
    -1554.29577636719, 
    -1601.76806640625, 
    -1646.88635253906, 
    -1684.98400878906, 
    -1696.66223144531, 
    -1672.51989746094, 
    -1718.88977050781, 
    -1813.208984375, 
    -1961.46215820312, 
    -1904.04992675781, 
    -1894.65417480469, 
    -1897.47583007812, 
    -1888.62976074219, 
    -1830.93273925781, 
    -1711.72302246094, 
    -1734.53552246094, 
    -1680.74450683594, 
    -1704.22009277344, 
    -1599.14819335938, 
    -1480.46423339844, 
    -1453.88220214844, 
    -1403.30786132812, 
    -1281.42651367188, 
    -1171.98132324219, 
    -1123.435546875, 
    -1008.06829833984, 
    -925.882446289062, 
    -933.773986816406, 
    -875.874877929688, 
    -769.886352539062, 
    -722.438415527344, 
    -589.721740722656, 
    -493.005920410156, 
    -459.493011474609, 
    -400.307037353516, 
    -406.000152587891, 
    -427.207733154297, 
    -409.547393798828, 
    -365.987335205078, 
    -312.313842773438, 
    -303.414184570312, 
    -334.39501953125, 
    -302.865325927734, 
    -265.353088378906, 
    -234.153350830078, 
    -294.365783691406, 
    -313.751739501953, 
    -86.7795028686523, 
    534.311096191406, 
    1048.29443359375, 
    987.738891601562, 
    1300.13891601562, 
    1032.36669921875, 
    1415.02770996094, 
    1881.77783203125, 
    1203.04443359375, 
    621.358093261719, 
    -540.769836425781, 
    -426.565521240234, 
    -318.508026123047, 
    -307.5595703125, 
    10.1116638183594, 
    302.436096191406, 
    433.347229003906, 
    850.291625976562, 
    727.288879394531, 
    642.566650390625, 
    -181.598007202148, 
    -2.41383028030396, 
    252.45556640625, 
    321.739532470703, 
    383.410552978516, 
    -57.5974273681641, 
    -290.127655029297, 
    660.747192382812, 
    614.180541992188, 
    652.91943359375, 
    224.720352172852, 
    -8.31170749664307, 
    807.927795410156, 
    844.516662597656, 
    577.725036621094, 
    341.711120605469, 
    142.519897460938, 
    -365.670684814453, 
    -51.403980255127, 
    236.152770996094, 
    113.55517578125, 
    -116.130905151367, 
    -303.889801025391, 
    -100.102973937988, 
    91.983772277832, 
    -70.0398788452148, 
    -178.538070678711, 
    -207.095489501953, 
    -175.496826171875, 
    -203.575393676758, 
    -153.374389648438, 
    -196.684692382812, 
    -324.677001953125, 
    -399.040405273438, 
    -290.024963378906, 
    -219.844390869141, 
    -82.9268341064453, 
    -80.899528503418, 
    -141.027633666992, 
    -78.6955947875977, 
    -99.0032119750977, 
    -120.856086730957, 
    -120.668922424316, 
    -231.563613891602, 
    -277.702178955078, 
    -197.637191772461, 
    -119.06761932373, 
    -165.742340087891, 
    -183.85920715332, 
    -153.784927368164, 
    -93.5536041259766, 
    -73.2145843505859, 
    -444.296875, 
    -1528.7607421875, 
    -2857.54858398438, 
    -3101.05029296875, 
    -3474.16186523438, 
    -3838.861328125, 
    -3873.9130859375, 
    -2569.70922851562, 
    -2458.91088867188, 
    -3201.9873046875, 
    -2456.412109375, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1619.05895996094, 
    -1492.37805175781, 
    -1453.77551269531, 
    -1348.86950683594, 
    -1429.99035644531, 
    -1550.91662597656, 
    -1655.53039550781, 
    -1712.25341796875, 
    -1738.90417480469, 
    -1644.88806152344, 
    -1623.96838378906, 
    -1747.43005371094, 
    -1806.61474609375, 
    -1823.63171386719, 
    -1831.3017578125, 
    -1820.38330078125, 
    -1794.66760253906, 
    -1705.12121582031, 
    -1677.98046875, 
    -1586.20092773438, 
    -1511.52502441406, 
    -1410.82995605469, 
    -1312.39709472656, 
    -1244.75402832031, 
    -1030.94274902344, 
    -1008.03540039062, 
    -899.626770019531, 
    -782.050354003906, 
    -551.192138671875, 
    -536.527282714844, 
    -596.913208007812, 
    -585.808288574219, 
    -560.930908203125, 
    -583.581970214844, 
    -632.952209472656, 
    -494.012115478516, 
    -504.260101318359, 
    -499.72509765625, 
    -539.308471679688, 
    -536.042907714844, 
    -571.683837890625, 
    -597.024963378906, 
    -357.289489746094, 
    -326.406646728516, 
    -381.204803466797, 
    -362.601715087891, 
    -304.531677246094, 
    -314.452850341797, 
    -285.3330078125, 
    -196.933471679688, 
    -86.3537750244141, 
    37.4585762023926, 
    424.419067382812, 
    505.661102294922, 
    784.450012207031, 
    1452.23608398438, 
    1590.59448242188, 
    1493.822265625, 
    885.734558105469, 
    -498.934661865234, 
    -285.692199707031, 
    -32.1931686401367, 
    150.599990844727, 
    142.58610534668, 
    388.516662597656, 
    840.561096191406, 
    554.91943359375, 
    248.125, 
    310.430541992188, 
    -371.588653564453, 
    634.663879394531, 
    178.566207885742, 
    45.7958679199219, 
    241.622222900391, 
    -91.7850494384766, 
    -349.231201171875, 
    -70.3430023193359, 
    180.441299438477, 
    602.383361816406, 
    689.536071777344, 
    18.4399375915527, 
    721.763854980469, 
    192.915481567383, 
    512.119445800781, 
    96.0741271972656, 
    -68.2988128662109, 
    -289.217864990234, 
    5.69866561889648, 
    -55.4869003295898, 
    -216.118835449219, 
    -329.610046386719, 
    -58.3026809692383, 
    -66.0104217529297, 
    -111.939933776855, 
    -171.864379882812, 
    -265.104705810547, 
    -249.205810546875, 
    -185.812149047852, 
    -169.473937988281, 
    -212.989105224609, 
    -294.587524414062, 
    -334.614013671875, 
    -395.360504150391, 
    -456.317657470703, 
    -249.72900390625, 
    -212.097259521484, 
    -142.109436035156, 
    -108.169563293457, 
    -192.089691162109, 
    -115.520286560059, 
    -160.546142578125, 
    -233.153106689453, 
    -259.726593017578, 
    -220.160949707031, 
    -214.478897094727, 
    -116.832572937012, 
    -157.523880004883, 
    -225.087615966797, 
    -251.285995483398, 
    -204.97346496582, 
    -245.768096923828, 
    -1107.0244140625, 
    -1840.10168457031, 
    -2987.63110351562, 
    -3374.67211914062, 
    -3459.75927734375, 
    -3924.67236328125, 
    -2936.75122070312, 
    -1893.89624023438, 
    -2684.39282226562, 
    -2325.0576171875, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1353.96655273438, 
    -1371.69982910156, 
    -1545.55798339844, 
    -1462.43103027344, 
    -1541.86645507812, 
    -1448.24182128906, 
    -1496.02856445312, 
    -1554.71081542969, 
    -1663.615234375, 
    -1681.31469726562, 
    -1620.52600097656, 
    -1622.04833984375, 
    -1628.94995117188, 
    -1594.22131347656, 
    -1547.96618652344, 
    -1717.89196777344, 
    -1745.05834960938, 
    -1705.64392089844, 
    -1599.91931152344, 
    -1502.06262207031, 
    -1354.31860351562, 
    -1191.56896972656, 
    -1024.66186523438, 
    -905.224365234375, 
    -763.739624023438, 
    -660.258117675781, 
    -438.555633544922, 
    -371.417419433594, 
    -301.338500976562, 
    -328.272705078125, 
    -359.510833740234, 
    -375.004577636719, 
    -367.028594970703, 
    -449.532836914062, 
    -595.8701171875, 
    -575.795104980469, 
    -561.98388671875, 
    -597.209777832031, 
    -631.299743652344, 
    -690.223999023438, 
    -761.946166992188, 
    -739.443908691406, 
    -666.586486816406, 
    -649.536193847656, 
    -726.988098144531, 
    -508.323944091797, 
    -364.418701171875, 
    -293.334045410156, 
    -276.176300048828, 
    -286.759918212891, 
    -185.406997680664, 
    -185.297210693359, 
    356.944885253906, 
    960.344421386719, 
    910.525024414062, 
    1312.42224121094, 
    1373.6416015625, 
    17.1430339813232, 
    -430.775787353516, 
    -104.486610412598, 
    188.202774047852, 
    348.783325195312, 
    330.186096191406, 
    427.424987792969, 
    492.911102294922, 
    382.516662597656, 
    -10.2483930587769, 
    211.038970947266, 
    -254.884948730469, 
    235.493179321289, 
    362.428955078125, 
    -148.87663269043, 
    -74.0898742675781, 
    -230.672271728516, 
    0.795822143554688, 
    -312.926208496094, 
    87.7671279907227, 
    228.063888549805, 
    429.299652099609, 
    -195.950042724609, 
    -151.552108764648, 
    303.819458007812, 
    452.511108398438, 
    64.0475463867188, 
    -222.492980957031, 
    -149.021697998047, 
    64.9761047363281, 
    31.7092056274414, 
    -281.06640625, 
    -462.847198486328, 
    -284.482269287109, 
    -249.549194335938, 
    -233.97053527832, 
    -349.900939941406, 
    -303.341888427734, 
    -202.098403930664, 
    -159.121673583984, 
    -214.630966186523, 
    -244.676742553711, 
    -293.831024169922, 
    -313.20703125, 
    -352.544128417969, 
    -405.282836914062, 
    -285.483612060547, 
    -219.321624755859, 
    -175.173492431641, 
    -189.902053833008, 
    -204.091918945312, 
    -318.277648925781, 
    -211.367492675781, 
    -298.994934082031, 
    -168.969116210938, 
    -186.863754272461, 
    -202.913986206055, 
    -200.934173583984, 
    -193.878631591797, 
    -231.334808349609, 
    -229.293121337891, 
    -268.965240478516, 
    -331.196624755859, 
    -2056.94482421875, 
    -2640.20581054688, 
    -3334.2978515625, 
    -3403.69458007812, 
    -3374.09448242188, 
    -3124.31298828125, 
    -2100.98022460938, 
    -1789.50329589844, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1039.5556640625, 
    -1081.43212890625, 
    -1251.3857421875, 
    -1438.86669921875, 
    -1487.00671386719, 
    -1410.06127929688, 
    -1531.09545898438, 
    -1482.49462890625, 
    -1553.30187988281, 
    -1596.88757324219, 
    -1600.56567382812, 
    -1529.70263671875, 
    -1437.42565917969, 
    -1390.09631347656, 
    -1291.28991699219, 
    -1304.98498535156, 
    -1366.57177734375, 
    -1496.23937988281, 
    -1460.10583496094, 
    -1283.25927734375, 
    -1122.25036621094, 
    -883.671325683594, 
    -687.512939453125, 
    -591.505554199219, 
    -380.280609130859, 
    -273.964385986328, 
    -234.010467529297, 
    -210.502365112305, 
    -192.624755859375, 
    -200.6298828125, 
    -200.492370605469, 
    -236.531616210938, 
    -260.1611328125, 
    -441.877624511719, 
    -592.955261230469, 
    -682.957336425781, 
    -700.414916992188, 
    -758.147888183594, 
    -867.476135253906, 
    -1007.96136474609, 
    -1004.65734863281, 
    -1182.90344238281, 
    -1155.43469238281, 
    -1286.83642578125, 
    -1120.61755371094, 
    -1045.73278808594, 
    -478.173767089844, 
    -387.343841552734, 
    -239.67399597168, 
    -334.189544677734, 
    -234.609085083008, 
    -171.855926513672, 
    87.1160888671875, 
    664.691650390625, 
    706.236083984375, 
    1237.86669921875, 
    -216.541412353516, 
    -397.308044433594, 
    109.590850830078, 
    506.483306884766, 
    549.011108398438, 
    487.311126708984, 
    401.175018310547, 
    182.042572021484, 
    -50.7891540527344, 
    268.228088378906, 
    -309.478790283203, 
    -416.462341308594, 
    -161.040588378906, 
    -211.171783447266, 
    -205.630462646484, 
    -262.951019287109, 
    -219.142913818359, 
    -132.372604370117, 
    -372.265045166016, 
    -206.97119140625, 
    -93.8735427856445, 
    -106.77840423584, 
    -200.591567993164, 
    -307.700866699219, 
    -41.9244422912598, 
    15.8033332824707, 
    266.641662597656, 
    -204.08464050293, 
    -192.730895996094, 
    55.048210144043, 
    24.2354373931885, 
    -320.913909912109, 
    -375.263916015625, 
    -146.077713012695, 
    -86.9619598388672, 
    -129.119552612305, 
    -284.238250732422, 
    -265.924865722656, 
    -207.981430053711, 
    -219.064224243164, 
    -189.497299194336, 
    -210.585678100586, 
    -299.142852783203, 
    -279.949249267578, 
    -349.391479492188, 
    -360.896636962891, 
    -299.280609130859, 
    -220.877532958984, 
    -171.765579223633, 
    -184.114669799805, 
    -182.071228027344, 
    -334.532409667969, 
    -237.384002685547, 
    -232.642517089844, 
    -183.051727294922, 
    -186.623962402344, 
    -198.892166137695, 
    -207.100799560547, 
    -198.368774414062, 
    -203.355438232422, 
    -417.670593261719, 
    -792.835205078125, 
    -2081.64892578125, 
    -2922.20043945312, 
    -2874.56640625, 
    -3644.57470703125, 
    -3810.39501953125, 
    -3045.40014648438, 
    -2779.14916992188, 
    -2345.55932617188, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2263.361328125, 
    -870.413208007812, 
    -792.835693359375, 
    -944.724853515625, 
    -1129.56469726562, 
    -1396.67321777344, 
    -1516.96557617188, 
    -1499.10656738281, 
    -1463.24560546875, 
    -1391.40161132812, 
    -1445.37365722656, 
    -1444.72644042969, 
    -1496.81225585938, 
    -1407.93115234375, 
    -1378.52490234375, 
    -1271.61486816406, 
    -1234.37915039062, 
    -1208.77661132812, 
    -1188.55041503906, 
    -1115.97839355469, 
    -968.86962890625, 
    -607.128479003906, 
    -405.581604003906, 
    -355.089599609375, 
    -315.760040283203, 
    -212.288452148438, 
    -180.557952880859, 
    -166.464874267578, 
    -152.53288269043, 
    -144.992782592773, 
    -152.006973266602, 
    -208.277709960938, 
    -197.524322509766, 
    -180.400833129883, 
    -287.285278320312, 
    -560.631408691406, 
    -774.264831542969, 
    -934.46044921875, 
    -1101.95776367188, 
    -1234.4541015625, 
    -1294.62561035156, 
    -1418.07727050781, 
    -1450.099609375, 
    -1464.16748046875, 
    -1414.84948730469, 
    -1343.0146484375, 
    -1195.08312988281, 
    -912.324096679688, 
    -261.509490966797, 
    -321.576416015625, 
    -239.272399902344, 
    -219.712051391602, 
    -243.402328491211, 
    -83.8315124511719, 
    357.989929199219, 
    694.269470214844, 
    247.890029907227, 
    -427.446899414062, 
    41.0160484313965, 
    273.364044189453, 
    117.142959594727, 
    432.702789306641, 
    550.099975585938, 
    494.016662597656, 
    30.4731273651123, 
    -253.431243896484, 
    -405.422760009766, 
    -382.281524658203, 
    -197.507843017578, 
    -222.800872802734, 
    -335.114105224609, 
    -266.336181640625, 
    -202.647506713867, 
    -198.714462280273, 
    -410.301055908203, 
    -258.429229736328, 
    -160.038864135742, 
    -181.383148193359, 
    -193.34260559082, 
    -242.063690185547, 
    -187.120513916016, 
    -161.853286743164, 
    -176.630187988281, 
    -248.441741943359, 
    -258.262817382812, 
    44.1934700012207, 
    -221.765029907227, 
    -325.256622314453, 
    -224.889938354492, 
    -160.904373168945, 
    -113.623985290527, 
    -180.196075439453, 
    -291.526763916016, 
    -282.855194091797, 
    -223.123687744141, 
    -235.664779663086, 
    -225.951263427734, 
    -237.258743286133, 
    -266.792572021484, 
    -271.967224121094, 
    -310.988220214844, 
    -322.287628173828, 
    -243.766342163086, 
    -171.951370239258, 
    -172.541854858398, 
    -196.942794799805, 
    -207.766784667969, 
    -259.486541748047, 
    -303.763977050781, 
    -245.119430541992, 
    -152.262969970703, 
    -187.188629150391, 
    -254.908630371094, 
    -280.648620605469, 
    -174.221527099609, 
    -294.382598876953, 
    -1115.35583496094, 
    -1647.29846191406, 
    -2567.16772460938, 
    -3176.19287109375, 
    -3426.87646484375, 
    -4285.1669921875, 
    -2894.98510742188, 
    -2987.77587890625, 
    -2373.53344726562, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2153.90966796875, 
    -1105.37707519531, 
    -905.234985351562, 
    -868.308959960938, 
    -902.038024902344, 
    -1042.76159667969, 
    -1324.32800292969, 
    -1510.83190917969, 
    -1439.76501464844, 
    -1393.28564453125, 
    -1408.51818847656, 
    -1379.16882324219, 
    -1360.99084472656, 
    -1371.27319335938, 
    -1353.08032226562, 
    -1308.89318847656, 
    -1215.88342285156, 
    -1107.38598632812, 
    -914.481628417969, 
    -501.066528320312, 
    -346.904388427734, 
    -327.167755126953, 
    -300.394378662109, 
    -289.516235351562, 
    -230.288925170898, 
    -188.210693359375, 
    -169.524963378906, 
    -139.600402832031, 
    -128.240737915039, 
    -112.10131072998, 
    -192.157043457031, 
    -133.20573425293, 
    -137.319961547852, 
    -148.766616821289, 
    -204.366363525391, 
    -403.388488769531, 
    -628.7548828125, 
    -779.015319824219, 
    -1013.88983154297, 
    -1086.83996582031, 
    -1086.67041015625, 
    -1318.76770019531, 
    -1452.18664550781, 
    -1454.30737304688, 
    -1434.17407226562, 
    -1434.966796875, 
    -1288.99133300781, 
    -608.659484863281, 
    -354.702789306641, 
    -414.421813964844, 
    -265.104339599609, 
    -209.777542114258, 
    -180.436126708984, 
    -123.829261779785, 
    -88.6021118164062, 
    555.069213867188, 
    -564.579528808594, 
    -306.588409423828, 
    525.386108398438, 
    644.980529785156, 
    431.658782958984, 
    -95.1747741699219, 
    -194.78205871582, 
    -207.477325439453, 
    -263.31396484375, 
    -299.776794433594, 
    -417.686126708984, 
    -207.778961181641, 
    -248.581100463867, 
    -280.260009765625, 
    -189.240905761719, 
    -233.375213623047, 
    -194.96435546875, 
    -423.958251953125, 
    -269.976348876953, 
    -176.23405456543, 
    -196.20588684082, 
    -218.634185791016, 
    -248.922424316406, 
    -188.971862792969, 
    -198.195465087891, 
    -225.350051879883, 
    -266.950714111328, 
    -345.282348632812, 
    -322.797027587891, 
    -301.21142578125, 
    -229.495162963867, 
    -155.260345458984, 
    -181.19841003418, 
    -148.357269287109, 
    -225.902679443359, 
    -300.591033935547, 
    -269.843231201172, 
    -209.302108764648, 
    -233.37825012207, 
    -201.433456420898, 
    -227.949798583984, 
    -265.363250732422, 
    -261.251281738281, 
    -264.266510009766, 
    -180.980346679688, 
    -205.476257324219, 
    -214.571105957031, 
    -186.181503295898, 
    -201.463241577148, 
    -247.491363525391, 
    -255.241897583008, 
    -242.939636230469, 
    -200.020401000977, 
    -201.724731445312, 
    -191.2578125, 
    -413.855072021484, 
    -389.993194580078, 
    -314.285064697266, 
    -1085.85681152344, 
    -1712.28820800781, 
    -2183.01733398438, 
    -2767.97924804688, 
    -3571.98022460938, 
    -4088.51318359375, 
    -2972.76416015625, 
    -3151.27172851562, 
    -2313.71044921875, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2065.86596679688, 
    -1256.23559570312, 
    -1013.92510986328, 
    -829.430786132812, 
    -789.888488769531, 
    -818.014038085938, 
    -908.779296875, 
    -1331.85278320312, 
    -1471.40710449219, 
    -1484.34326171875, 
    -1340.71447753906, 
    -1408.83642578125, 
    -1237.43249511719, 
    -1314.49780273438, 
    -1271.10998535156, 
    -1133.35107421875, 
    -923.780334472656, 
    -620.503051757812, 
    -282.0126953125, 
    -292.924896240234, 
    -330.308959960938, 
    -328.032257080078, 
    -288.210235595703, 
    -228.228530883789, 
    -189.798034667969, 
    -155.661819458008, 
    -130.83447265625, 
    -107.127281188965, 
    -88.448112487793, 
    -91.9393463134766, 
    -105.713966369629, 
    -123.327613830566, 
    -99.0445098876953, 
    -112.242050170898, 
    -110.455749511719, 
    -163.503326416016, 
    -277.889343261719, 
    -629.103515625, 
    -730.0673828125, 
    -865.55615234375, 
    -988.458557128906, 
    -1154.4951171875, 
    -1355.13842773438, 
    -1414.69067382812, 
    -1463.18200683594, 
    -1440.1572265625, 
    -1432.48950195312, 
    -1389.24157714844, 
    -1188.72290039062, 
    -658.759887695312, 
    -283.079315185547, 
    -279.340942382812, 
    -313.464599609375, 
    -431.690460205078, 
    -402.404327392578, 
    -424.483673095703, 
    -406.696960449219, 
    289.523132324219, 
    -144.194946289062, 
    -267.735443115234, 
    -274.433074951172, 
    -284.608612060547, 
    -264.846008300781, 
    -246.312225341797, 
    -251.530319213867, 
    -322.870513916016, 
    -246.654678344727, 
    -264.939666748047, 
    -260.255981445312, 
    -258.265472412109, 
    -234.576370239258, 
    -225.58186340332, 
    -370.34130859375, 
    -230.430648803711, 
    -218.409790039062, 
    -265.034423828125, 
    -268.027191162109, 
    -249.376617431641, 
    -186.561569213867, 
    -198.317886352539, 
    -237.834899902344, 
    -303.998291015625, 
    -348.747375488281, 
    -299.707092285156, 
    -226.936904907227, 
    -150.456420898438, 
    -178.72834777832, 
    -203.272171020508, 
    -175.619003295898, 
    -293.708465576172, 
    -305.96484375, 
    -217.269775390625, 
    -205.766189575195, 
    -213.607391357422, 
    -208.22966003418, 
    -255.514663696289, 
    -286.684265136719, 
    -247.115325927734, 
    -257.524261474609, 
    -280.727111816406, 
    -236.641754150391, 
    -234.065170288086, 
    -206.194381713867, 
    -199.974380493164, 
    -228.464965820312, 
    -235.031280517578, 
    -191.551406860352, 
    -206.16259765625, 
    -265.310638427734, 
    -274.524688720703, 
    -587.953735351562, 
    -808.191650390625, 
    -1327.2431640625, 
    -1786.87097167969, 
    -2174.77978515625, 
    -2493.27905273438, 
    -2843.87670898438, 
    -3215.81127929688, 
    -2744.6279296875, 
    -3026.72778320312, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1636.45703125, 
    -1381.80212402344, 
    -1276.80834960938, 
    -953.402465820312, 
    -821.770690917969, 
    -789.358154296875, 
    -760.751586914062, 
    -834.141479492188, 
    -1085.408203125, 
    -1355.09338378906, 
    -1412.03198242188, 
    -1254.84753417969, 
    -1281.80651855469, 
    -1189.67163085938, 
    -991.282531738281, 
    -589.264831542969, 
    -376.619750976562, 
    -307.766387939453, 
    -226.100128173828, 
    -291.180908203125, 
    -291.167694091797, 
    -271.736968994141, 
    -215.181533813477, 
    -178.377883911133, 
    -143.495529174805, 
    -116.933815002441, 
    -82.7237014770508, 
    -64.8662261962891, 
    -58.7799263000488, 
    -61.3405265808105, 
    -88.2800216674805, 
    -78.1071548461914, 
    -96.3492050170898, 
    -107.669990539551, 
    -174.589752197266, 
    -172.152038574219, 
    -244.110275268555, 
    -395.737701416016, 
    -566.35400390625, 
    -731.663635253906, 
    -896.468872070312, 
    -1112.53894042969, 
    -1239.37463378906, 
    -1343.1533203125, 
    -1415.94445800781, 
    -1464.76721191406, 
    -1494.09558105469, 
    -1338.25427246094, 
    -526.60986328125, 
    -368.635284423828, 
    -358.364410400391, 
    -408.524200439453, 
    -445.929016113281, 
    -491.319244384766, 
    -580.550109863281, 
    -486.517059326172, 
    -308.9814453125, 
    -263.669738769531, 
    -286.493103027344, 
    -313.764495849609, 
    -383.277435302734, 
    -298.345062255859, 
    -258.933532714844, 
    -268.842712402344, 
    -315.675018310547, 
    -235.330749511719, 
    -249.566299438477, 
    -263.851470947266, 
    -261.855407714844, 
    -253.331466674805, 
    -296.33544921875, 
    -392.967895507812, 
    -287.09814453125, 
    -202.401138305664, 
    -227.734375, 
    -265.436859130859, 
    -234.570907592773, 
    -222.879028320312, 
    -221.546524047852, 
    -258.252624511719, 
    -300.071990966797, 
    -292.780975341797, 
    -228.209075927734, 
    -159.47917175293, 
    -154.139373779297, 
    -202.416732788086, 
    -206.004852294922, 
    -184.910293579102, 
    -293.401184082031, 
    -297.542358398438, 
    -192.377212524414, 
    -216.321685791016, 
    -210.889663696289, 
    -291.256286621094, 
    -282.715545654297, 
    -324.923767089844, 
    -448.182434082031, 
    -416.420623779297, 
    -310.097717285156, 
    -267.463470458984, 
    -248.15869140625, 
    -215.126831054688, 
    -221.741714477539, 
    -255.546417236328, 
    -200.393417358398, 
    -218.243835449219, 
    -241.532669067383, 
    -369.111053466797, 
    -590.710144042969, 
    -1322.66772460938, 
    -1678.64611816406, 
    -1874.58471679688, 
    -2218.91333007812, 
    -2471.68383789062, 
    -2688.3525390625, 
    -2771.56591796875, 
    -2330.8466796875, 
    -2437.27490234375, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -1363.92687988281, 
    -1358.93249511719, 
    -1365.29943847656, 
    -1107.11511230469, 
    -861.81005859375, 
    -832.393798828125, 
    -641.65576171875, 
    -678.33984375, 
    -796.59130859375, 
    -928.266357421875, 
    -1278.89245605469, 
    -1307.30651855469, 
    -1131.06970214844, 
    -826.850769042969, 
    -338.431213378906, 
    -306.248260498047, 
    -373.335479736328, 
    -251.00764465332, 
    -219.233291625977, 
    -257.886260986328, 
    -245.578384399414, 
    -246.872512817383, 
    -201.888061523438, 
    -148.853286743164, 
    -97.1578674316406, 
    -77.4829177856445, 
    -53.7613906860352, 
    -7.94443798065186, 
    -38.6915588378906, 
    -41.1147918701172, 
    -46.3032150268555, 
    -84.3723449707031, 
    -159.207626342773, 
    -113.503433227539, 
    -183.030578613281, 
    -234.3046875, 
    -267.647766113281, 
    -407.089416503906, 
    -471.283905029297, 
    -672.232788085938, 
    -881.028503417969, 
    -1082.72485351562, 
    -1196.49597167969, 
    -1276.28698730469, 
    -1367.57409667969, 
    -1449.79174804688, 
    -1377.33459472656, 
    -701.968078613281, 
    -383.523193359375, 
    -401.609375, 
    -424.888732910156, 
    -418.300262451172, 
    -432.800659179688, 
    -406.888275146484, 
    -333.60791015625, 
    -300.940460205078, 
    -262.891967773438, 
    -280.377899169922, 
    -318.854858398438, 
    -405.406036376953, 
    -409.585723876953, 
    -282.917419433594, 
    -296.665435791016, 
    -348.951599121094, 
    -290.767822265625, 
    -261.066589355469, 
    -264.675659179688, 
    -254.128295898438, 
    -262.890777587891, 
    -296.422912597656, 
    -348.468170166016, 
    -292.171142578125, 
    -255.558319091797, 
    -270.635528564453, 
    -286.477233886719, 
    -232.742630004883, 
    -234.434158325195, 
    -202.629913330078, 
    -283.114715576172, 
    -300.878692626953, 
    -254.683990478516, 
    -188.508316040039, 
    -159.390319824219, 
    -186.666000366211, 
    -192.266677856445, 
    -233.709213256836, 
    -217.607940673828, 
    -298.708953857422, 
    -334.650970458984, 
    -233.907485961914, 
    -174.935577392578, 
    -242.309158325195, 
    -317.729553222656, 
    -309.466522216797, 
    -359.639587402344, 
    -482.180786132812, 
    -388.957458496094, 
    -242.78776550293, 
    -211.258743286133, 
    -227.148193359375, 
    -223.206893920898, 
    -172.432113647461, 
    -271.030609130859, 
    -269.246673583984, 
    -292.833801269531, 
    -306.005462646484, 
    -466.151336669922, 
    -1330.93518066406, 
    -1785.72302246094, 
    -1994.42456054688, 
    -2173.8662109375, 
    -2466.1591796875, 
    -2675.63671875, 
    -2683.78491210938, 
    -2634.26440429688, 
    -2368.77221679688, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300,
  
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2250.68383789062, 
    -1400.50634765625, 
    -1424.14929199219, 
    -1321.79235839844, 
    -1278.04321289062, 
    -951.636901855469, 
    -731.353088378906, 
    -722.617004394531, 
    -655.805480957031, 
    -663.283325195312, 
    -745.808044433594, 
    -931.327575683594, 
    -933.998413085938, 
    -638.528076171875, 
    -309.360107421875, 
    -319.787231445312, 
    -417.896453857422, 
    -322.08056640625, 
    -211.88020324707, 
    -200.595336914062, 
    -189.751861572266, 
    -244.622039794922, 
    -274.150268554688, 
    -199.157623291016, 
    -95.0760116577148, 
    -85.334602355957, 
    -49.0030174255371, 
    -0.100000001490116, 
    -2.00420618057251, 
    -5.57215213775635, 
    -2.94372344017029, 
    -95.0428619384766, 
    -80.348991394043, 
    -74.1234588623047, 
    -124.209915161133, 
    -228.062225341797, 
    -247.419845581055, 
    -342.585418701172, 
    -480.039184570312, 
    -623.585388183594, 
    -737.005798339844, 
    -832.127197265625, 
    -938.916259765625, 
    -1024.86022949219, 
    -1195.23474121094, 
    -1379.82934570312, 
    -1432.76391601562, 
    -999.169860839844, 
    -387.697631835938, 
    -408.95263671875, 
    -393.076080322266, 
    -333.392852783203, 
    -320.229827880859, 
    -304.96875, 
    -296.968017578125, 
    -293.372894287109, 
    -276.126281738281, 
    -304.462280273438, 
    -650.504455566406, 
    -817.973815917969, 
    -568.504028320312, 
    -572.588928222656, 
    -546.495361328125, 
    -563.104431152344, 
    -411.15380859375, 
    -491.656524658203, 
    -542.475402832031, 
    -407.462799072266, 
    -266.425140380859, 
    -273.710510253906, 
    -347.135070800781, 
    -290.478820800781, 
    -321.451995849609, 
    -586.927307128906, 
    -298.601501464844, 
    -410.456787109375, 
    -539.658569335938, 
    -481.442993164062, 
    -283.261047363281, 
    -293.221466064453, 
    -171.817077636719, 
    -196.205322265625, 
    -187.550796508789, 
    -200.877670288086, 
    -195.607086181641, 
    -223.419052124023, 
    -191.009490966797, 
    -277.759063720703, 
    -377.121459960938, 
    -253.715957641602, 
    -241.039123535156, 
    -303.030914306641, 
    -303.614776611328, 
    -306.833587646484, 
    -318.075164794922, 
    -380.322265625, 
    -329.408599853516, 
    -269.145233154297, 
    -191.028244018555, 
    -267.344665527344, 
    -295.507598876953, 
    -211.538146972656, 
    -333.675506591797, 
    -321.088409423828, 
    -353.575286865234, 
    -416.252746582031, 
    -1075.7607421875, 
    -1741.50634765625, 
    -2209.19897460938, 
    -2288.50415039062, 
    -2362.89868164062, 
    -2504.26513671875, 
    -2709.0634765625, 
    -2768.16186523438, 
    -2323.65698242188, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300, 
    -2300 ;
}
