// Sample Icebin parameter file.  Place in [rundir]/config/icebin.cdl
//

netcdf icebin {
variables:
    // Setup methods (in ectl) to be run after symlinks are
    // created and before ModelE is launched.
    // Names of these attributes can be whatever you like
    int setups ;
        setups:landice = "ectl.xsetup.pism_landice.xsetup";

    // ModelE-specific variables cover all ice sheets
    int m.info ;

        // Determines mapping between GCM's elevation classes,
        // and the elevation classes that are passed to IceBin.
        //
        // legacy [1]: A single elevation class for ice not associated
        //             with elevation classes.
        // sealand[2]: Two elevation classes, providing separation
        //             between ocean and land portions of an atmosphere
        //             grid cell.
        // ec[n]:      A set of IceBin-defined elevation classes
        m.info:segments = "legacy,sealand,ec";

        m.info:grid = "input-file:landice/pismsheet_g20_icebin_in.nc";

        // Where IceBin may write stuff
        m.info:output_dir = "output-dir:icebin";

        // Set to "f" and IceBin will pass a zero SMB and
        // appropriately zero B.C. to the ice sheet.  This is for
        // testing.
        m.info:use_smb = "t" ;

    // Additional variables agument m.greenland.info from main icebin_in
    // These variables are specific to Greenland
    int m.greenland.info ;
        // Output for greenland-specific stuff
        m.greenland.info:output_dir = "output-dir:greenland";

        // The ice model with which we are coupling.
        // See IceCoupler::Type [DISMAL, PISM, ISSM, WRITER]
        m.greenland.info:ice_coupler = "PISM" ;

        // Should we upate the elevation field in update_ice_sheet()?
        // Normally, yes.  But in some TEST CASES ONLY --- when the SMB
        // field was created with a different set of elevations than the
        // ice model is using --- then this can cause problems in the
        // generated SMB fields.
        // See IceModel_PISM::update_elevation
        m.greenland.info:update_elevation = "f" ;

        // Variable currently in icebin_in, but maybe they should be moved here.
        // m.greenland.info:interp_grid = "EXCH" ;
        // m.greenland.info:interp_style = "Z_INTERP" ;
        // Also: hcdefs, indexingHC

    // Variables specific to the ModelE side of the coupling
    double m.greenland.modele ;

        // Should ModelE prepare for Dirichlet or Neumann boundary
        // conditions with the dynamic ice model?
        // See 
        m.greenland.modele:coupling_type = "DIRICHLET_BC" ;

    double m.greenland.pism ;
        // Command-line arguments provided to PISM upon initialization
        // Paths will be resolved for filenames in this list.
        m.greenland.pism:i = "input-file:pism/std-greenland/g20km_10ka.nc" ;
        m.greenland.pism:skip = "" ;
        m.greenland.pism:skip_max = "10" ;
        m.greenland.pism:surface = "given" ;
        m.greenland.pism:surface_given_file = "input-file:pism/std-greenland/pism_Greenland_5km_v1.1.nc" ;
        m.greenland.pism:calving = "ocean_kill" ;
        m.greenland.pism:ocean_kill_file = "input-file:pism/std-greenland/pism_Greenland_5km_v1.1.nc" ;
        m.greenland.pism:sia_e = "3.0" ;
        m.greenland.pism:ts_file = "output-file:greenland/ts_g20km_10ka_run2.nc" ;
        m.greenland.pism:ts_times = "0:1:1000" ;
        m.greenland.pism:extra_file = "output-file:greenland/ex_g20km_10ka_run2.nc" ;
        m.greenland.pism:extra_times = "0:.1:1000" ;
        m.greenland.pism:extra_vars = "climatic_mass_balance,ice_surface_temp,diffusivity,temppabase,tempicethk_basal,bmelt,tillwat,csurf,mask,thk,topg,usurf" ;
        m.greenland.pism:o = "g20km_10ka_run2.nc" ;
    double m.greenland.dismal ;
        m.greenland.dismal:output_dir = "dismal_out2" ;

}
